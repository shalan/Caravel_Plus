magic
tech sky130A
magscale 1 2
timestamp 1610138030
<< nwell >>
rect 0 616613 352 617179
rect 0 615525 352 616091
rect 0 614437 352 615003
rect 0 613349 352 613915
rect 0 612261 352 612827
rect 0 611173 352 611739
rect 0 610085 352 610651
rect 0 608997 352 609563
rect 0 607909 352 608475
rect 0 606821 352 607387
rect 0 605733 352 606299
rect 0 604645 352 605211
rect 0 603878 352 604123
rect 0 603802 6608 603878
rect 0 603557 5136 603802
rect 0 602790 352 603035
rect 0 602714 78920 602790
rect 0 602469 10380 602714
rect 0 601381 352 601947
rect 0 600293 352 600859
rect 0 599205 352 599771
rect 0 598117 352 598683
rect 0 597350 352 597595
rect 0 597029 2836 597350
rect 0 595941 352 596507
rect 0 594853 352 595419
rect 0 593765 352 594331
rect 0 592677 352 593243
rect 0 591589 352 592155
rect 0 590501 352 591067
rect 0 589413 352 589979
rect 0 588325 352 588891
rect 0 587237 352 587803
rect 0 586149 352 586715
rect 0 585617 513 585627
rect 0 585382 1824 585617
rect 0 585306 6608 585382
rect 0 585061 352 585306
rect 0 583973 352 584539
rect 0 582885 352 583451
rect 0 581797 352 582363
rect 0 581030 1824 581275
rect 0 580954 50400 581030
rect 0 580709 352 580954
rect 0 579621 352 580187
rect 0 578854 1824 579099
rect 0 578778 46260 578854
rect 0 578543 3940 578778
rect 0 578533 513 578543
rect 0 577766 1824 578011
rect 0 577690 47640 577766
rect 0 577445 352 577690
rect 0 576357 352 576923
rect 0 575269 352 575835
rect 0 574181 352 574747
rect 0 573093 352 573659
rect 0 572005 352 572571
rect 0 570917 352 571483
rect 0 569829 352 570395
rect 0 568741 352 569307
rect 0 567653 352 568219
rect 0 566886 2008 567131
rect 0 566810 42672 566886
rect 0 566565 4124 566810
rect 0 565477 352 566043
rect 0 564389 352 564955
rect 0 563301 352 563867
rect 0 562213 352 562779
rect 0 561125 352 561691
rect 0 560037 352 560603
rect 0 558949 352 559515
rect 0 558182 352 558427
rect 0 558106 2100 558182
rect 0 557871 2008 558106
rect 0 557861 513 557871
rect 0 556773 352 557339
rect 0 555685 352 556251
rect 0 554597 352 555163
rect 0 553509 352 554075
rect 0 552421 352 552987
rect 0 551333 352 551899
rect 0 550245 352 550811
rect 0 549157 352 549723
rect 0 548390 2836 548635
rect 0 548314 54540 548390
rect 0 548069 5412 548314
rect 0 547302 1180 547547
rect 0 547226 6240 547302
rect 0 546991 5596 547226
rect 0 546981 513 546991
rect 0 545893 352 546459
rect 0 545126 352 545371
rect 0 545050 22432 545126
rect 0 544805 3204 545050
rect 0 544038 2008 544283
rect 0 543962 3112 544038
rect 0 543717 352 543962
rect 0 542629 352 543195
rect 0 541541 352 542107
rect 0 540453 352 541019
rect 0 539365 352 539931
rect 0 538277 352 538843
rect 0 537189 352 537755
rect 0 536101 352 536667
rect 0 535013 352 535579
rect 0 533925 352 534491
rect 0 532837 352 533403
rect 0 531749 352 532315
rect 0 530661 352 531227
rect 0 529573 352 530139
rect 0 528806 1824 529051
rect 0 528730 2744 528806
rect 0 528485 352 528730
rect 0 527397 352 527963
rect 0 526865 513 526875
rect 0 526630 8448 526865
rect 0 526554 20868 526630
rect 0 526309 352 526554
rect 0 525542 1824 525787
rect 0 525466 14060 525542
rect 0 525221 3020 525466
rect 0 524133 352 524699
rect 0 523366 2008 523611
rect 0 523290 25100 523366
rect 0 523045 352 523290
rect 0 522202 2836 522523
rect 0 521957 352 522202
rect 0 521190 1824 521435
rect 0 521114 24824 521190
rect 0 520869 352 521114
rect 0 519781 352 520347
rect 0 518693 352 519259
rect 0 517605 352 518171
rect 0 516838 352 517083
rect 0 516527 1824 516838
rect 0 516517 513 516527
rect 0 515750 352 515995
rect 0 515674 89684 515750
rect 0 515429 5320 515674
rect 0 514341 352 514907
rect 0 513253 352 513819
rect 0 512165 352 512731
rect 0 511077 352 511643
rect 0 510310 352 510555
rect 0 510234 19488 510310
rect 0 509999 5596 510234
rect 0 509989 1985 509999
rect 0 508901 352 509467
rect 0 508134 352 508379
rect 0 508058 13416 508134
rect 0 507813 1824 508058
rect 0 506725 352 507291
rect 0 505637 352 506203
rect 0 504549 2836 505115
rect 0 503461 352 504027
rect 0 502694 2008 502939
rect 0 502618 47088 502694
rect 0 502383 2100 502618
rect 0 502373 513 502383
rect 0 501606 3020 501851
rect 0 501530 33656 501606
rect 0 501285 2836 501530
rect 0 500197 352 500763
rect 0 499430 352 499675
rect 0 499354 5964 499430
rect 0 499109 3296 499354
rect 0 498342 2836 498587
rect 0 498266 8816 498342
rect 0 498021 352 498266
rect 0 497254 2008 497499
rect 0 497178 15624 497254
rect 0 496933 352 497178
rect 0 496166 1824 496411
rect 0 496090 22064 496166
rect 0 495845 352 496090
rect 0 495313 513 495323
rect 0 495078 2836 495313
rect 0 495002 3848 495078
rect 0 494757 1180 495002
rect 0 493990 352 494235
rect 0 493914 113236 493990
rect 0 493679 3112 493914
rect 0 493669 1985 493679
rect 0 492902 1824 493147
rect 0 492826 9460 492902
rect 0 492581 352 492826
rect 0 491493 352 492059
rect 0 490726 352 490971
rect 0 490650 15716 490726
rect 0 490415 1824 490650
rect 0 490405 513 490415
rect 0 489317 352 489883
rect 0 488229 352 488795
rect 0 487141 352 487707
rect 0 486053 352 486619
rect 0 484965 352 485531
rect 0 483877 352 484443
rect 0 483345 513 483355
rect 0 483110 1824 483345
rect 0 483034 11116 483110
rect 0 482789 352 483034
rect 0 482022 3848 482267
rect 0 481946 11208 482022
rect 0 481701 352 481946
rect 0 480934 2008 481179
rect 0 480858 56012 480934
rect 0 480613 5596 480858
rect 0 479846 2836 480091
rect 0 479770 28044 479846
rect 0 479525 352 479770
rect 0 478993 513 479003
rect 0 478758 1824 478993
rect 0 478682 22616 478758
rect 0 478437 352 478682
rect 0 477670 8448 477915
rect 0 477594 11024 477670
rect 0 477349 352 477594
rect 0 476261 352 476827
rect 0 475173 352 475739
rect 0 474406 352 474651
rect 0 474085 3480 474406
rect 0 473318 352 473563
rect 0 473242 8448 473318
rect 0 472997 5596 473242
rect 0 472465 513 472475
rect 0 472230 5504 472465
rect 0 472154 11576 472230
rect 0 471909 352 472154
rect 0 471142 352 471387
rect 0 470821 2836 471142
rect 0 470054 2836 470299
rect 0 469978 15072 470054
rect 0 469733 2652 469978
rect 0 468645 352 469211
rect 0 467557 352 468123
rect 0 466469 352 467035
rect 0 465381 352 465947
rect 0 464293 352 464859
rect 0 463205 352 463771
rect 0 462117 352 462683
rect 0 461029 352 461595
rect 0 459941 352 460507
rect 0 459174 3204 459419
rect 0 459098 55460 459174
rect 0 458853 352 459098
rect 0 458321 513 458331
rect 0 458086 4492 458321
rect 0 458010 70548 458086
rect 0 457765 352 458010
rect 0 456677 352 457243
rect 0 455589 352 456155
rect 0 454822 352 455067
rect 0 454501 3664 454822
rect 0 453734 2836 453979
rect 0 453658 22340 453734
rect 0 453413 352 453658
rect 0 452325 352 452891
rect 0 451558 2836 451803
rect 0 451482 16820 451558
rect 0 451237 352 451482
rect 0 450470 352 450715
rect 0 450394 42120 450470
rect 0 450159 2008 450394
rect 0 450149 513 450159
rect 0 449382 352 449627
rect 0 449306 19396 449382
rect 0 449071 2100 449306
rect 0 449061 513 449071
rect 0 447973 352 448539
rect 0 446885 352 447451
rect 0 446118 1824 446363
rect 0 446042 42580 446118
rect 0 445797 352 446042
rect 0 444709 352 445275
rect 0 443621 352 444187
rect 0 442533 352 443099
rect 0 441445 352 442011
rect 0 440678 352 440923
rect 0 440602 6884 440678
rect 0 440357 1824 440602
rect 0 439269 352 439835
rect 0 438181 352 438747
rect 0 437649 513 437659
rect 0 437414 1824 437649
rect 0 437338 5596 437414
rect 0 437093 352 437338
rect 0 436005 352 436571
rect 0 434917 352 435483
rect 0 433829 352 434395
rect 0 433062 352 433307
rect 0 432986 36416 433062
rect 0 432741 3480 432986
rect 0 431653 352 432219
rect 0 431121 513 431131
rect 0 430886 1824 431121
rect 0 430810 3940 430886
rect 0 430565 352 430810
rect 0 429798 352 430043
rect 0 429722 12864 429798
rect 0 429487 5596 429722
rect 0 429477 2997 429487
rect 0 428945 513 428955
rect 0 428710 1824 428945
rect 0 428634 66500 428710
rect 0 428389 352 428634
rect 0 427301 352 427867
rect 0 426534 352 426779
rect 0 426458 8448 426534
rect 0 426213 2008 426458
rect 0 425446 352 425691
rect 0 425370 6148 425446
rect 0 425125 3664 425370
rect 0 424037 352 424603
rect 0 422949 352 423515
rect 0 421861 352 422427
rect 0 420773 352 421339
rect 0 420006 2468 420251
rect 0 419930 5872 420006
rect 0 419685 352 419930
rect 0 419153 513 419163
rect 0 418842 1824 419153
rect 0 418597 352 418842
rect 0 417509 352 418075
rect 0 416666 3204 416987
rect 0 416421 2192 416666
rect 0 415333 352 415899
rect 0 414490 2836 414811
rect 0 414245 352 414490
rect 0 413157 2836 413723
rect 0 412069 352 412635
rect 0 410981 352 411547
rect 0 409893 352 410459
rect 0 408805 352 409371
rect 0 407717 352 408283
rect 0 406629 352 407195
rect 0 405541 352 406107
rect 0 404453 352 405019
rect 0 403365 352 403931
rect 0 402277 352 402843
rect 0 401189 352 401755
rect 0 400422 352 400667
rect 0 400346 10104 400422
rect 0 400111 3940 400346
rect 0 400101 513 400111
rect 0 399013 352 399579
rect 0 397925 352 398491
rect 0 396837 352 397403
rect 0 395749 352 396315
rect 0 394661 352 395227
rect 0 393573 352 394139
rect 0 392485 352 393051
rect 0 391397 352 391963
rect 0 390309 352 390875
rect 0 389221 352 389787
rect 0 388133 352 388699
rect 0 387366 1824 387611
rect 0 387290 92628 387366
rect 0 387045 352 387290
rect 0 385957 352 386523
rect 0 385425 513 385435
rect 0 385190 1824 385425
rect 0 385114 50032 385190
rect 0 384869 352 385114
rect 0 383781 352 384347
rect 0 382693 352 383259
rect 0 381605 352 382171
rect 0 380838 352 381083
rect 0 380762 31264 380838
rect 0 380527 4768 380762
rect 0 380517 513 380527
rect 0 379429 352 379995
rect 0 378662 352 378907
rect 0 378586 16360 378662
rect 0 378341 3664 378586
rect 0 377574 2008 377819
rect 0 377498 11576 377574
rect 0 377253 352 377498
rect 0 376165 352 376731
rect 0 375077 352 375643
rect 0 373989 352 374555
rect 0 372901 352 373467
rect 0 371813 352 372379
rect 0 370725 352 371291
rect 0 369637 352 370203
rect 0 368549 352 369115
rect 0 367461 352 368027
rect 0 366373 352 366939
rect 0 365285 352 365851
rect 0 364197 352 364763
rect 0 363109 352 363675
rect 0 362021 352 362587
rect 0 360933 352 361499
rect 0 359845 352 360411
rect 0 358757 352 359323
rect 0 357669 352 358235
rect 0 356581 352 357147
rect 0 355493 352 356059
rect 0 354405 352 354971
rect 0 353317 352 353883
rect 0 352229 352 352795
rect 0 351141 352 351707
rect 0 350053 352 350619
rect 0 348965 352 349531
rect 0 347877 352 348443
rect 0 346789 352 347355
rect 0 345701 352 346267
rect 0 344613 352 345179
rect 0 343525 352 344091
rect 0 342437 352 343003
rect 0 341349 352 341915
rect 0 340261 352 340827
rect 0 339173 352 339739
rect 0 338085 352 338651
rect 0 336997 352 337563
rect 0 335909 352 336475
rect 0 334821 352 335387
rect 0 333733 352 334299
rect 0 332645 352 333211
rect 0 331557 352 332123
rect 0 330469 352 331035
rect 0 329381 352 329947
rect 0 328293 352 328859
rect 0 327205 352 327771
rect 0 326117 352 326683
rect 0 325029 352 325595
rect 0 323941 352 324507
rect 0 322853 352 323419
rect 0 321765 352 322331
rect 0 320677 352 321243
rect 0 319589 352 320155
rect 0 318501 352 319067
rect 0 317413 352 317979
rect 0 316325 352 316891
rect 0 315237 352 315803
rect 0 314149 352 314715
rect 0 313061 352 313627
rect 0 311973 352 312539
rect 0 310885 352 311451
rect 0 309797 352 310363
rect 0 308709 352 309275
rect 0 307621 352 308187
rect 0 306533 352 307099
rect 0 305445 352 306011
rect 0 304357 352 304923
rect 0 303269 352 303835
rect 0 302181 352 302747
rect 0 301093 352 301659
rect 0 300005 352 300571
rect 0 298917 352 299483
rect 0 297829 352 298395
rect 0 296741 352 297307
rect 0 295653 352 296219
rect 0 294565 352 295131
rect 0 293477 352 294043
rect 0 292389 352 292955
rect 0 291301 352 291867
rect 0 290213 352 290779
rect 0 289446 2836 289691
rect 0 289370 16636 289446
rect 0 289125 352 289370
rect 0 288037 352 288603
rect 0 286949 352 287515
rect 0 285861 352 286427
rect 0 284773 352 285339
rect 0 283685 352 284251
rect 0 282597 352 283163
rect 0 281509 352 282075
rect 0 280421 352 280987
rect 0 279333 352 279899
rect 0 278245 352 278811
rect 0 277157 352 277723
rect 0 276069 352 276635
rect 0 274981 352 275547
rect 0 273893 352 274459
rect 0 272805 352 273371
rect 0 271717 352 272283
rect 0 270629 352 271195
rect 0 269541 352 270107
rect 0 268453 352 269019
rect 0 267365 352 267931
rect 0 266277 352 266843
rect 0 265189 352 265755
rect 0 264101 352 264667
rect 0 263013 352 263579
rect 0 261925 352 262491
rect 0 260837 352 261403
rect 0 259749 352 260315
rect 0 258661 352 259227
rect 0 257573 352 258139
rect 0 256485 352 257051
rect 0 255397 352 255963
rect 0 254309 352 254875
rect 0 253221 352 253787
rect 0 252133 352 252699
rect 0 251045 352 251611
rect 0 249957 352 250523
rect 0 248869 352 249435
rect 0 247781 352 248347
rect 0 246693 352 247259
rect 0 245605 352 246171
rect 0 244517 352 245083
rect 0 243429 352 243995
rect 0 242341 352 242907
rect 0 241253 352 241819
rect 0 240165 352 240731
rect 0 239077 352 239643
rect 0 237989 352 238555
rect 0 236901 352 237467
rect 0 235813 352 236379
rect 0 234725 352 235291
rect 0 233637 352 234203
rect 0 232549 352 233115
rect 0 231461 352 232027
rect 0 230373 352 230939
rect 0 229285 352 229851
rect 0 228197 352 228763
rect 0 227109 352 227675
rect 0 226021 352 226587
rect 0 224933 352 225499
rect 0 223845 352 224411
rect 0 222757 352 223323
rect 0 221669 352 222235
rect 0 220581 352 221147
rect 0 219493 352 220059
rect 0 218405 352 218971
rect 0 217317 352 217883
rect 0 216229 352 216795
rect 0 215141 352 215707
rect 0 214053 352 214619
rect 0 212965 352 213531
rect 0 211877 352 212443
rect 0 210789 352 211355
rect 0 209701 352 210267
rect 0 208613 352 209179
rect 0 207525 352 208091
rect 0 206437 352 207003
rect 0 205349 352 205915
rect 0 204261 352 204827
rect 0 203173 352 203739
rect 0 202085 352 202651
rect 0 200997 352 201563
rect 0 199909 352 200475
rect 0 198821 352 199387
rect 0 197733 352 198299
rect 0 196645 352 197211
rect 0 195557 352 196123
rect 0 194469 352 195035
rect 0 193381 352 193947
rect 0 192293 352 192859
rect 0 191205 352 191771
rect 0 190117 352 190683
rect 0 189029 352 189595
rect 0 187941 352 188507
rect 0 186853 352 187419
rect 0 185765 352 186331
rect 0 184677 352 185243
rect 0 183589 352 184155
rect 0 182501 352 183067
rect 0 181413 352 181979
rect 0 180646 352 180891
rect 0 180325 2192 180646
rect 0 179558 1824 179803
rect 0 179482 3112 179558
rect 0 179237 352 179482
rect 0 178470 1824 178715
rect 0 178394 5780 178470
rect 0 178149 352 178394
rect 0 177382 2836 177627
rect 0 177306 3296 177382
rect 0 177061 352 177306
rect 0 175973 352 176539
rect 0 175206 352 175451
rect 0 175130 8264 175206
rect 0 174895 1824 175130
rect 0 174885 513 174895
rect 0 174118 352 174363
rect 0 174042 5228 174118
rect 0 173797 2652 174042
rect 0 172709 352 173275
rect 0 171942 352 172187
rect 0 171866 15072 171942
rect 0 171631 1824 171866
rect 0 171621 513 171631
rect 0 170854 352 171099
rect 0 170778 33564 170854
rect 0 170533 4124 170778
rect 0 169445 352 170011
rect 0 168357 352 168923
rect 0 167269 352 167835
rect 0 166502 352 166747
rect 0 166426 24640 166502
rect 0 166191 3756 166426
rect 0 166181 513 166191
rect 0 165414 352 165659
rect 0 165338 3848 165414
rect 0 165093 3480 165338
rect 0 164005 352 164571
rect 0 163473 513 163483
rect 0 163238 1824 163473
rect 0 163162 3848 163238
rect 0 162917 352 163162
rect 0 161829 352 162395
rect 0 161062 352 161307
rect 0 160741 2008 161062
rect 0 159974 2836 160219
rect 0 159898 3020 159974
rect 0 159653 352 159898
rect 0 158565 352 159131
rect 0 157477 352 158043
rect 0 156710 1824 156955
rect 0 156634 16820 156710
rect 0 156399 2008 156634
rect 0 156389 513 156399
rect 0 155301 352 155867
rect 0 154213 352 154779
rect 0 153125 352 153691
rect 0 152037 352 152603
rect 0 151270 352 151515
rect 0 151194 95388 151270
rect 0 150959 5596 151194
rect 0 150949 513 150959
rect 0 149871 2008 150427
rect 0 149861 513 149871
rect 0 148773 352 149339
rect 0 147685 3204 148251
rect 0 146918 2652 147163
rect 0 146842 53620 146918
rect 0 146597 352 146842
rect 0 145830 352 146075
rect 0 145754 3848 145830
rect 0 145509 3664 145754
rect 0 144742 352 144987
rect 0 144666 35680 144742
rect 0 144421 5596 144666
rect 0 143654 352 143899
rect 0 143578 36140 143654
rect 0 143343 8264 143578
rect 0 143333 513 143343
rect 0 142566 352 142811
rect 0 142490 47456 142566
rect 0 142255 1824 142490
rect 0 142245 513 142255
rect 0 141157 352 141723
rect 0 140069 352 140635
rect 0 138981 352 139547
rect 0 138214 2836 138459
rect 0 138138 14520 138214
rect 0 137893 3480 138138
rect 0 137126 352 137371
rect 0 137050 25100 137126
rect 0 136805 2008 137050
rect 0 136038 2836 136283
rect 0 135962 25284 136038
rect 0 135717 352 135962
rect 0 134950 2836 135195
rect 0 134874 70180 134950
rect 0 134629 352 134874
rect 0 133862 352 134107
rect 0 133786 33380 133862
rect 0 133541 1824 133786
rect 0 132774 2836 133019
rect 0 132698 4768 132774
rect 0 132453 352 132698
rect 0 131686 2836 131931
rect 0 131365 4768 131686
rect 0 130598 2836 130843
rect 0 130522 8356 130598
rect 0 130277 2192 130522
rect 0 129510 2836 129755
rect 0 129434 8264 129510
rect 0 129189 352 129434
rect 0 128422 2836 128667
rect 0 128346 16820 128422
rect 0 128101 352 128346
rect 0 127334 2836 127579
rect 0 127258 14244 127334
rect 0 127013 352 127258
rect 0 126246 352 126491
rect 0 126170 21052 126246
rect 0 125935 3296 126170
rect 0 125925 513 125935
rect 0 124837 352 125403
rect 0 123749 352 124315
rect 0 122982 2836 123227
rect 0 122906 50216 122982
rect 0 122671 5136 122906
rect 0 122661 1985 122671
rect 0 121894 352 122139
rect 0 121573 4124 121894
rect 0 120485 352 121051
rect 0 119397 352 119963
rect 0 118309 352 118875
rect 0 117221 352 117787
rect 0 116133 352 116699
rect 0 115045 352 115611
rect 0 113957 352 114523
rect 0 112869 352 113435
rect 0 111781 352 112347
rect 0 110693 352 111259
rect 0 109605 352 110171
rect 0 108517 352 109083
rect 0 107429 352 107995
rect 0 106341 352 106907
rect 0 105253 352 105819
rect 0 104165 352 104731
rect 0 103077 352 103643
rect 0 101989 352 102555
rect 0 100901 352 101467
rect 0 99813 352 100379
rect 0 98725 352 99291
rect 0 97637 352 98203
rect 0 96549 352 97115
rect 0 95461 352 96027
rect 0 94373 352 94939
rect 0 93285 352 93851
rect 0 92197 352 92763
rect 0 91109 352 91675
rect 0 90021 352 90587
rect 0 88933 352 89499
rect 0 87845 352 88411
rect 0 86757 352 87323
rect 0 85669 352 86235
rect 0 84581 352 85147
rect 0 83493 352 84059
rect 0 82405 352 82971
rect 0 81317 352 81883
rect 0 80229 352 80795
rect 0 79141 352 79707
rect 0 78053 352 78619
rect 0 76965 352 77531
rect 0 75877 352 76443
rect 0 74789 352 75355
rect 0 73701 352 74267
rect 0 72613 352 73179
rect 0 71525 352 72091
rect 0 70437 352 71003
rect 0 69349 352 69915
rect 0 68261 352 68827
rect 0 67173 352 67739
rect 0 66085 352 66651
rect 0 64997 352 65563
rect 0 63909 352 64475
rect 0 62821 352 63387
rect 0 61733 352 62299
rect 0 60645 352 61211
rect 0 59557 352 60123
rect 0 58469 352 59035
rect 0 57381 352 57947
rect 0 56293 352 56859
rect 0 55205 352 55771
rect 0 54117 352 54683
rect 0 53029 352 53595
rect 0 51941 352 52507
rect 0 50853 352 51419
rect 0 49765 352 50331
rect 0 48677 352 49243
rect 0 47589 352 48155
rect 0 46501 352 47067
rect 0 45413 352 45979
rect 0 44325 352 44891
rect 0 43237 352 43803
rect 0 42149 352 42715
rect 0 41061 352 41627
rect 0 39973 352 40539
rect 0 38885 352 39451
rect 0 37797 352 38363
rect 0 36709 352 37275
rect 0 35621 352 36187
rect 0 34533 352 35099
rect 0 33445 352 34011
rect 0 32357 352 32923
rect 0 31269 352 31835
rect 0 30181 352 30747
rect 0 29093 352 29659
rect 0 28005 352 28571
rect 0 26917 352 27483
rect 0 25829 352 26395
rect 0 24741 352 25307
rect 0 23653 352 24219
rect 0 22565 352 23131
rect 0 21477 352 22043
rect 0 20389 352 20955
rect 0 19301 352 19867
rect 0 18213 352 18779
rect 0 17125 352 17691
rect 0 16037 352 16603
rect 0 14949 352 15515
rect 0 13861 352 14427
rect 0 12773 352 13339
rect 0 11685 352 12251
rect 0 10597 352 11163
rect 0 9509 352 10075
rect 0 8421 352 8987
rect 0 7333 352 7899
rect 0 6245 352 6811
rect 0 5157 352 5723
rect 0 4069 352 4635
rect 0 2981 352 3547
rect 0 2138 352 2459
<< obsli1 >>
rect 38 1989 577953 617559
<< obsm1 >>
rect 38 892 577965 617568
<< metal2 >>
rect 2356 0 2412 800
rect 9256 0 9312 800
rect 16248 0 16304 800
rect 23240 0 23296 800
rect 30232 0 30288 800
rect 37224 0 37280 800
rect 44216 0 44272 800
rect 51208 0 51264 800
rect 58200 0 58256 800
rect 65192 0 65248 800
rect 72184 0 72240 800
rect 79176 0 79232 800
rect 86168 0 86224 800
rect 93160 0 93216 800
rect 100152 0 100208 800
rect 107144 0 107200 800
rect 114136 0 114192 800
rect 121128 0 121184 800
rect 128120 0 128176 800
rect 135112 0 135168 800
rect 142104 0 142160 800
rect 149004 0 149060 800
rect 155996 0 156052 800
rect 162988 0 163044 800
rect 169980 0 170036 800
rect 176972 0 177028 800
rect 183964 0 184020 800
rect 190956 0 191012 800
rect 197948 0 198004 800
rect 204940 0 204996 800
rect 211932 0 211988 800
rect 218924 0 218980 800
rect 225916 0 225972 800
rect 232908 0 232964 800
rect 239900 0 239956 800
rect 246892 0 246948 800
rect 253884 0 253940 800
rect 260876 0 260932 800
rect 267868 0 267924 800
rect 274860 0 274916 800
rect 281852 0 281908 800
rect 288844 0 288900 800
rect 295744 0 295800 800
rect 302736 0 302792 800
rect 309728 0 309784 800
rect 316720 0 316776 800
rect 323712 0 323768 800
rect 330704 0 330760 800
rect 337696 0 337752 800
rect 344688 0 344744 800
rect 351680 0 351736 800
rect 358672 0 358728 800
rect 365664 0 365720 800
rect 372656 0 372712 800
rect 379648 0 379704 800
rect 386640 0 386696 800
rect 393632 0 393688 800
rect 400624 0 400680 800
rect 407616 0 407672 800
rect 414608 0 414664 800
rect 421600 0 421656 800
rect 428592 0 428648 800
rect 435584 0 435640 800
rect 442484 0 442540 800
rect 449476 0 449532 800
rect 456468 0 456524 800
rect 463460 0 463516 800
rect 470452 0 470508 800
rect 477444 0 477500 800
rect 484436 0 484492 800
rect 491428 0 491484 800
rect 498420 0 498476 800
rect 505412 0 505468 800
rect 512404 0 512460 800
rect 519396 0 519452 800
rect 526388 0 526444 800
rect 533380 0 533436 800
rect 540372 0 540428 800
rect 547364 0 547420 800
rect 554356 0 554412 800
rect 561348 0 561404 800
rect 568340 0 568396 800
rect 575332 0 575388 800
<< obsm2 >>
rect 334 856 577778 617574
rect 334 800 2300 856
rect 2468 800 9200 856
rect 9368 800 16192 856
rect 16360 800 23184 856
rect 23352 800 30176 856
rect 30344 800 37168 856
rect 37336 800 44160 856
rect 44328 800 51152 856
rect 51320 800 58144 856
rect 58312 800 65136 856
rect 65304 800 72128 856
rect 72296 800 79120 856
rect 79288 800 86112 856
rect 86280 800 93104 856
rect 93272 800 100096 856
rect 100264 800 107088 856
rect 107256 800 114080 856
rect 114248 800 121072 856
rect 121240 800 128064 856
rect 128232 800 135056 856
rect 135224 800 142048 856
rect 142216 800 148948 856
rect 149116 800 155940 856
rect 156108 800 162932 856
rect 163100 800 169924 856
rect 170092 800 176916 856
rect 177084 800 183908 856
rect 184076 800 190900 856
rect 191068 800 197892 856
rect 198060 800 204884 856
rect 205052 800 211876 856
rect 212044 800 218868 856
rect 219036 800 225860 856
rect 226028 800 232852 856
rect 233020 800 239844 856
rect 240012 800 246836 856
rect 247004 800 253828 856
rect 253996 800 260820 856
rect 260988 800 267812 856
rect 267980 800 274804 856
rect 274972 800 281796 856
rect 281964 800 288788 856
rect 288956 800 295688 856
rect 295856 800 302680 856
rect 302848 800 309672 856
rect 309840 800 316664 856
rect 316832 800 323656 856
rect 323824 800 330648 856
rect 330816 800 337640 856
rect 337808 800 344632 856
rect 344800 800 351624 856
rect 351792 800 358616 856
rect 358784 800 365608 856
rect 365776 800 372600 856
rect 372768 800 379592 856
rect 379760 800 386584 856
rect 386752 800 393576 856
rect 393744 800 400568 856
rect 400736 800 407560 856
rect 407728 800 414552 856
rect 414720 800 421544 856
rect 421712 800 428536 856
rect 428704 800 435528 856
rect 435696 800 442428 856
rect 442596 800 449420 856
rect 449588 800 456412 856
rect 456580 800 463404 856
rect 463572 800 470396 856
rect 470564 800 477388 856
rect 477556 800 484380 856
rect 484548 800 491372 856
rect 491540 800 498364 856
rect 498532 800 505356 856
rect 505524 800 512348 856
rect 512516 800 519340 856
rect 519508 800 526332 856
rect 526500 800 533324 856
rect 533492 800 540316 856
rect 540484 800 547308 856
rect 547476 800 554300 856
rect 554468 800 561292 856
rect 561460 800 568284 856
rect 568452 800 575276 856
rect 575444 800 577778 856
<< obsm3 >>
rect 511 851 577601 617473
<< metal4 >>
rect 3142 2128 3462 617488
rect 18502 2128 18822 617488
rect 33862 2128 34182 617488
rect 49222 2128 49542 617488
rect 64582 2128 64902 617488
rect 79942 2128 80262 617488
rect 95302 2128 95622 617488
rect 110662 2128 110982 617488
rect 126022 2128 126342 617488
rect 141382 2128 141702 617488
rect 156742 2128 157062 617488
rect 172102 2128 172422 617488
rect 187462 2128 187782 617488
rect 202822 2128 203142 617488
rect 218182 2128 218502 617488
rect 233542 2128 233862 617488
rect 248902 2128 249222 617488
rect 264262 2128 264582 617488
rect 279622 2128 279942 617488
rect 294982 2128 295302 617488
rect 310342 2128 310662 617488
rect 325702 2128 326022 617488
rect 341062 2128 341382 617488
rect 356422 2128 356742 617488
rect 371782 2128 372102 617488
rect 387142 2128 387462 617488
rect 402502 2128 402822 617488
rect 417862 2128 418182 617488
rect 433222 2128 433542 617488
rect 448582 2128 448902 617488
rect 463942 2128 464262 617488
rect 479302 2128 479622 617488
rect 494662 2128 494982 617488
rect 510022 2128 510342 617488
rect 525382 2128 525702 617488
rect 540742 2128 541062 617488
rect 556102 2128 556422 617488
rect 571462 2128 571782 617488
<< obsm4 >>
rect 2489 2048 3062 616589
rect 3542 2048 18422 616589
rect 18902 2048 33782 616589
rect 34262 2048 49142 616589
rect 49622 2048 64502 616589
rect 64982 2048 79862 616589
rect 80342 2048 95222 616589
rect 95702 2048 110582 616589
rect 111062 2048 125942 616589
rect 126422 2048 141302 616589
rect 141782 2048 156662 616589
rect 157142 2048 172022 616589
rect 172502 2048 187382 616589
rect 187862 2048 202742 616589
rect 203222 2048 218102 616589
rect 218582 2048 233462 616589
rect 233942 2048 248822 616589
rect 249302 2048 264182 616589
rect 264662 2048 279542 616589
rect 280022 2048 294902 616589
rect 295382 2048 310262 616589
rect 310742 2048 325622 616589
rect 326102 2048 340982 616589
rect 341462 2048 356342 616589
rect 356822 2048 371702 616589
rect 372182 2048 387062 616589
rect 387542 2048 402422 616589
rect 402902 2048 417782 616589
rect 418262 2048 433142 616589
rect 433622 2048 448502 616589
rect 448982 2048 463862 616589
rect 464342 2048 479222 616589
rect 479702 2048 494582 616589
rect 495062 2048 509942 616589
rect 510422 2048 525302 616589
rect 525782 2048 540662 616589
rect 541142 2048 556022 616589
rect 556502 2048 571382 616589
rect 571862 2048 575163 616589
rect 2489 1939 575163 2048
<< labels >>
rlabel metal2 s 449476 0 449532 800 6 A[0]
port 1 nsew signal input
rlabel metal2 s 519396 0 519452 800 6 A[10]
port 2 nsew signal input
rlabel metal2 s 526388 0 526444 800 6 A[11]
port 3 nsew signal input
rlabel metal2 s 533380 0 533436 800 6 A[12]
port 4 nsew signal input
rlabel metal2 s 456468 0 456524 800 6 A[1]
port 5 nsew signal input
rlabel metal2 s 463460 0 463516 800 6 A[2]
port 6 nsew signal input
rlabel metal2 s 470452 0 470508 800 6 A[3]
port 7 nsew signal input
rlabel metal2 s 477444 0 477500 800 6 A[4]
port 8 nsew signal input
rlabel metal2 s 484436 0 484492 800 6 A[5]
port 9 nsew signal input
rlabel metal2 s 491428 0 491484 800 6 A[6]
port 10 nsew signal input
rlabel metal2 s 498420 0 498476 800 6 A[7]
port 11 nsew signal input
rlabel metal2 s 505412 0 505468 800 6 A[8]
port 12 nsew signal input
rlabel metal2 s 512404 0 512460 800 6 A[9]
port 13 nsew signal input
rlabel metal2 s 540372 0 540428 800 6 CLK
port 14 nsew signal input
rlabel metal2 s 225916 0 225972 800 6 Di[0]
port 15 nsew signal input
rlabel metal2 s 295744 0 295800 800 6 Di[10]
port 16 nsew signal input
rlabel metal2 s 302736 0 302792 800 6 Di[11]
port 17 nsew signal input
rlabel metal2 s 309728 0 309784 800 6 Di[12]
port 18 nsew signal input
rlabel metal2 s 316720 0 316776 800 6 Di[13]
port 19 nsew signal input
rlabel metal2 s 323712 0 323768 800 6 Di[14]
port 20 nsew signal input
rlabel metal2 s 330704 0 330760 800 6 Di[15]
port 21 nsew signal input
rlabel metal2 s 337696 0 337752 800 6 Di[16]
port 22 nsew signal input
rlabel metal2 s 344688 0 344744 800 6 Di[17]
port 23 nsew signal input
rlabel metal2 s 351680 0 351736 800 6 Di[18]
port 24 nsew signal input
rlabel metal2 s 358672 0 358728 800 6 Di[19]
port 25 nsew signal input
rlabel metal2 s 232908 0 232964 800 6 Di[1]
port 26 nsew signal input
rlabel metal2 s 365664 0 365720 800 6 Di[20]
port 27 nsew signal input
rlabel metal2 s 372656 0 372712 800 6 Di[21]
port 28 nsew signal input
rlabel metal2 s 379648 0 379704 800 6 Di[22]
port 29 nsew signal input
rlabel metal2 s 386640 0 386696 800 6 Di[23]
port 30 nsew signal input
rlabel metal2 s 393632 0 393688 800 6 Di[24]
port 31 nsew signal input
rlabel metal2 s 400624 0 400680 800 6 Di[25]
port 32 nsew signal input
rlabel metal2 s 407616 0 407672 800 6 Di[26]
port 33 nsew signal input
rlabel metal2 s 414608 0 414664 800 6 Di[27]
port 34 nsew signal input
rlabel metal2 s 421600 0 421656 800 6 Di[28]
port 35 nsew signal input
rlabel metal2 s 428592 0 428648 800 6 Di[29]
port 36 nsew signal input
rlabel metal2 s 239900 0 239956 800 6 Di[2]
port 37 nsew signal input
rlabel metal2 s 435584 0 435640 800 6 Di[30]
port 38 nsew signal input
rlabel metal2 s 442484 0 442540 800 6 Di[31]
port 39 nsew signal input
rlabel metal2 s 246892 0 246948 800 6 Di[3]
port 40 nsew signal input
rlabel metal2 s 253884 0 253940 800 6 Di[4]
port 41 nsew signal input
rlabel metal2 s 260876 0 260932 800 6 Di[5]
port 42 nsew signal input
rlabel metal2 s 267868 0 267924 800 6 Di[6]
port 43 nsew signal input
rlabel metal2 s 274860 0 274916 800 6 Di[7]
port 44 nsew signal input
rlabel metal2 s 281852 0 281908 800 6 Di[8]
port 45 nsew signal input
rlabel metal2 s 288844 0 288900 800 6 Di[9]
port 46 nsew signal input
rlabel metal2 s 2356 0 2412 800 6 Do[0]
port 47 nsew signal output
rlabel metal2 s 72184 0 72240 800 6 Do[10]
port 48 nsew signal output
rlabel metal2 s 79176 0 79232 800 6 Do[11]
port 49 nsew signal output
rlabel metal2 s 86168 0 86224 800 6 Do[12]
port 50 nsew signal output
rlabel metal2 s 93160 0 93216 800 6 Do[13]
port 51 nsew signal output
rlabel metal2 s 100152 0 100208 800 6 Do[14]
port 52 nsew signal output
rlabel metal2 s 107144 0 107200 800 6 Do[15]
port 53 nsew signal output
rlabel metal2 s 114136 0 114192 800 6 Do[16]
port 54 nsew signal output
rlabel metal2 s 121128 0 121184 800 6 Do[17]
port 55 nsew signal output
rlabel metal2 s 128120 0 128176 800 6 Do[18]
port 56 nsew signal output
rlabel metal2 s 135112 0 135168 800 6 Do[19]
port 57 nsew signal output
rlabel metal2 s 9256 0 9312 800 6 Do[1]
port 58 nsew signal output
rlabel metal2 s 142104 0 142160 800 6 Do[20]
port 59 nsew signal output
rlabel metal2 s 149004 0 149060 800 6 Do[21]
port 60 nsew signal output
rlabel metal2 s 155996 0 156052 800 6 Do[22]
port 61 nsew signal output
rlabel metal2 s 162988 0 163044 800 6 Do[23]
port 62 nsew signal output
rlabel metal2 s 169980 0 170036 800 6 Do[24]
port 63 nsew signal output
rlabel metal2 s 176972 0 177028 800 6 Do[25]
port 64 nsew signal output
rlabel metal2 s 183964 0 184020 800 6 Do[26]
port 65 nsew signal output
rlabel metal2 s 190956 0 191012 800 6 Do[27]
port 66 nsew signal output
rlabel metal2 s 197948 0 198004 800 6 Do[28]
port 67 nsew signal output
rlabel metal2 s 204940 0 204996 800 6 Do[29]
port 68 nsew signal output
rlabel metal2 s 16248 0 16304 800 6 Do[2]
port 69 nsew signal output
rlabel metal2 s 211932 0 211988 800 6 Do[30]
port 70 nsew signal output
rlabel metal2 s 218924 0 218980 800 6 Do[31]
port 71 nsew signal output
rlabel metal2 s 23240 0 23296 800 6 Do[3]
port 72 nsew signal output
rlabel metal2 s 30232 0 30288 800 6 Do[4]
port 73 nsew signal output
rlabel metal2 s 37224 0 37280 800 6 Do[5]
port 74 nsew signal output
rlabel metal2 s 44216 0 44272 800 6 Do[6]
port 75 nsew signal output
rlabel metal2 s 51208 0 51264 800 6 Do[7]
port 76 nsew signal output
rlabel metal2 s 58200 0 58256 800 6 Do[8]
port 77 nsew signal output
rlabel metal2 s 65192 0 65248 800 6 Do[9]
port 78 nsew signal output
rlabel metal2 s 575332 0 575388 800 6 EN
port 79 nsew signal input
rlabel metal2 s 547364 0 547420 800 6 WE[0]
port 80 nsew signal input
rlabel metal2 s 554356 0 554412 800 6 WE[1]
port 81 nsew signal input
rlabel metal2 s 561348 0 561404 800 6 WE[2]
port 82 nsew signal input
rlabel metal2 s 568340 0 568396 800 6 WE[3]
port 83 nsew signal input
rlabel metal4 s 556102 2128 556422 617488 6 VPWR
port 84 nsew power bidirectional
rlabel metal4 s 525382 2128 525702 617488 6 VPWR
port 85 nsew power bidirectional
rlabel metal4 s 494662 2128 494982 617488 6 VPWR
port 86 nsew power bidirectional
rlabel metal4 s 463942 2128 464262 617488 6 VPWR
port 87 nsew power bidirectional
rlabel metal4 s 433222 2128 433542 617488 6 VPWR
port 88 nsew power bidirectional
rlabel metal4 s 402502 2128 402822 617488 6 VPWR
port 89 nsew power bidirectional
rlabel metal4 s 371782 2128 372102 617488 6 VPWR
port 90 nsew power bidirectional
rlabel metal4 s 341062 2128 341382 617488 6 VPWR
port 91 nsew power bidirectional
rlabel metal4 s 310342 2128 310662 617488 6 VPWR
port 92 nsew power bidirectional
rlabel metal4 s 279622 2128 279942 617488 6 VPWR
port 93 nsew power bidirectional
rlabel metal4 s 248902 2128 249222 617488 6 VPWR
port 94 nsew power bidirectional
rlabel metal4 s 218182 2128 218502 617488 6 VPWR
port 95 nsew power bidirectional
rlabel metal4 s 187462 2128 187782 617488 6 VPWR
port 96 nsew power bidirectional
rlabel metal4 s 156742 2128 157062 617488 6 VPWR
port 97 nsew power bidirectional
rlabel metal4 s 126022 2128 126342 617488 6 VPWR
port 98 nsew power bidirectional
rlabel metal4 s 95302 2128 95622 617488 6 VPWR
port 99 nsew power bidirectional
rlabel metal4 s 64582 2128 64902 617488 6 VPWR
port 100 nsew power bidirectional
rlabel metal4 s 33862 2128 34182 617488 6 VPWR
port 101 nsew power bidirectional
rlabel metal4 s 3142 2128 3462 617488 6 VPWR
port 102 nsew power bidirectional
rlabel metal4 s 571462 2128 571782 617488 6 VGND
port 103 nsew ground bidirectional
rlabel metal4 s 540742 2128 541062 617488 6 VGND
port 104 nsew ground bidirectional
rlabel metal4 s 510022 2128 510342 617488 6 VGND
port 105 nsew ground bidirectional
rlabel metal4 s 479302 2128 479622 617488 6 VGND
port 106 nsew ground bidirectional
rlabel metal4 s 448582 2128 448902 617488 6 VGND
port 107 nsew ground bidirectional
rlabel metal4 s 417862 2128 418182 617488 6 VGND
port 108 nsew ground bidirectional
rlabel metal4 s 387142 2128 387462 617488 6 VGND
port 109 nsew ground bidirectional
rlabel metal4 s 356422 2128 356742 617488 6 VGND
port 110 nsew ground bidirectional
rlabel metal4 s 325702 2128 326022 617488 6 VGND
port 111 nsew ground bidirectional
rlabel metal4 s 294982 2128 295302 617488 6 VGND
port 112 nsew ground bidirectional
rlabel metal4 s 264262 2128 264582 617488 6 VGND
port 113 nsew ground bidirectional
rlabel metal4 s 233542 2128 233862 617488 6 VGND
port 114 nsew ground bidirectional
rlabel metal4 s 202822 2128 203142 617488 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 172102 2128 172422 617488 6 VGND
port 116 nsew ground bidirectional
rlabel metal4 s 141382 2128 141702 617488 6 VGND
port 117 nsew ground bidirectional
rlabel metal4 s 110662 2128 110982 617488 6 VGND
port 118 nsew ground bidirectional
rlabel metal4 s 79942 2128 80262 617488 6 VGND
port 119 nsew ground bidirectional
rlabel metal4 s 49222 2128 49542 617488 6 VGND
port 120 nsew ground bidirectional
rlabel metal4 s 18502 2128 18822 617488 6 VGND
port 121 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 577965 617574
string LEFview TRUE
string GDS_FILE ../gds/RAM_6Kx32.gds
string GDS_END 1274001762
string GDS_START 212328
<< end >>

