magic
tech sky130A
magscale 1 2
timestamp 1611017171
<< nwell >>
rect 0 616613 577836 617179
rect 0 615525 577836 616091
rect 0 614993 323065 615003
rect 0 614447 577836 614993
rect 0 614437 290497 614447
rect 0 613905 180833 613915
rect 0 613359 577836 613905
rect 0 613349 120021 613359
rect 0 612817 146241 612827
rect 0 612271 577836 612817
rect 0 612261 111097 612271
rect 0 611729 114041 611739
rect 0 611183 577836 611729
rect 0 611173 126093 611183
rect 0 610641 154705 610651
rect 0 610095 577836 610641
rect 0 610085 110545 610095
rect 0 609553 129405 609563
rect 0 609007 577836 609553
rect 0 608997 133453 609007
rect 0 608465 117629 608475
rect 0 607919 577836 608465
rect 0 607909 126553 607919
rect 0 607377 113857 607387
rect 0 606831 577836 607377
rect 0 606821 120573 606831
rect 0 606289 123609 606299
rect 0 605743 577836 606289
rect 0 605733 112569 605743
rect 0 605201 73929 605211
rect 0 604655 577836 605201
rect 0 604645 63901 604655
rect 0 604113 55621 604123
rect 0 603567 577836 604113
rect 0 603557 32437 603567
rect 0 603025 23513 603035
rect 0 602479 577836 603025
rect 0 602469 19925 602479
rect 0 601937 7413 601947
rect 0 601391 577836 601937
rect 0 601381 13945 601391
rect 0 600849 11185 600859
rect 0 600303 577836 600849
rect 0 600293 81565 600303
rect 0 599761 5849 599771
rect 0 599215 577836 599761
rect 0 599205 2353 599215
rect 0 598673 6033 598683
rect 0 598127 577836 598673
rect 0 598117 22777 598127
rect 0 597585 11553 597595
rect 0 597039 577836 597585
rect 0 597029 34277 597039
rect 0 596497 54241 596507
rect 0 595951 577836 596497
rect 0 595941 697 595951
rect 0 595409 7321 595419
rect 0 594863 577836 595409
rect 0 594853 19649 594863
rect 0 594321 29585 594331
rect 0 593775 577836 594321
rect 0 593765 56725 593775
rect 0 593233 1709 593243
rect 0 592687 577836 593233
rect 0 592677 13577 592687
rect 0 592145 76137 592155
rect 0 591599 577836 592145
rect 0 591589 513 591599
rect 0 591057 23421 591067
rect 0 590511 577836 591057
rect 0 590501 8701 590511
rect 0 589969 44857 589979
rect 0 589423 577836 589969
rect 0 589413 23145 589423
rect 0 588881 20017 588891
rect 0 588335 577836 588881
rect 0 588325 6309 588335
rect 0 587793 14497 587803
rect 0 587247 577836 587793
rect 0 587237 30873 587247
rect 0 586705 513 586715
rect 0 586159 577836 586705
rect 0 586149 17441 586159
rect 0 585617 54609 585627
rect 0 585071 577836 585617
rect 0 585061 789 585071
rect 0 584529 10449 584539
rect 0 583983 577836 584529
rect 0 583973 43845 583983
rect 0 583441 6953 583451
rect 0 582895 577836 583441
rect 0 582885 13669 582895
rect 0 582353 22133 582363
rect 0 581807 577836 582353
rect 0 581797 4193 581807
rect 0 581265 55897 581275
rect 0 580719 577836 581265
rect 0 580709 47249 580719
rect 0 580177 4929 580187
rect 0 579631 577836 580177
rect 0 579621 19281 579631
rect 0 579089 1801 579099
rect 0 578543 577836 579089
rect 0 578533 18085 578543
rect 0 578001 60773 578011
rect 0 577455 577836 578001
rect 0 577445 4285 577455
rect 0 576913 41085 576923
rect 0 576367 577836 576913
rect 0 576357 14221 576367
rect 0 575825 26273 575835
rect 0 575279 577836 575825
rect 0 575269 7781 575279
rect 0 574737 1249 574747
rect 0 574191 577836 574737
rect 0 574181 97297 574191
rect 0 573649 55621 573659
rect 0 573103 577836 573649
rect 0 573093 59301 573103
rect 0 572561 46697 572571
rect 0 572015 577836 572561
rect 0 572005 789 572015
rect 0 571473 15877 571483
rect 0 570927 577836 571473
rect 0 570917 84693 570927
rect 0 570385 14405 570395
rect 0 569839 577836 570385
rect 0 569829 1985 569839
rect 0 569297 7413 569307
rect 0 568751 577836 569297
rect 0 568741 4285 568751
rect 0 568209 10909 568219
rect 0 567663 577836 568209
rect 0 567653 7505 567663
rect 0 567121 60497 567131
rect 0 566575 577836 567121
rect 0 566565 25813 566575
rect 0 566033 513 566043
rect 0 565487 577836 566033
rect 0 565477 15417 565487
rect 0 564945 18085 564955
rect 0 564399 577836 564945
rect 0 564389 49273 564399
rect 0 563857 1801 563867
rect 0 563311 577836 563857
rect 0 563301 21397 563311
rect 0 562769 25813 562779
rect 0 562223 577836 562769
rect 0 562213 22961 562223
rect 0 561681 11093 561691
rect 0 561135 577836 561681
rect 0 561125 11829 561135
rect 0 560593 4101 560603
rect 0 560047 577836 560593
rect 0 560037 20569 560047
rect 0 559505 1433 559515
rect 0 558959 577836 559505
rect 0 558949 35565 558959
rect 0 558417 4653 558427
rect 0 557871 577836 558417
rect 0 557861 13393 557871
rect 0 557329 10357 557339
rect 0 556783 577836 557329
rect 0 556773 21397 556783
rect 0 556241 789 556251
rect 0 555695 577836 556241
rect 0 555685 7505 555695
rect 0 555153 35473 555163
rect 0 554607 577836 555153
rect 0 554597 55069 554607
rect 0 554065 23145 554075
rect 0 553519 577836 554065
rect 0 553509 65557 553519
rect 0 552977 1617 552987
rect 0 552431 577836 552977
rect 0 552421 4561 552431
rect 0 551889 72641 551899
rect 0 551343 577836 551889
rect 0 551333 15417 551343
rect 0 550801 21121 550811
rect 0 550255 577836 550801
rect 0 550245 4561 550255
rect 0 549713 26457 549723
rect 0 549167 577836 549713
rect 0 549157 8057 549167
rect 0 548625 7413 548635
rect 0 548079 577836 548625
rect 0 548069 973 548079
rect 0 547537 37497 547547
rect 0 546991 577836 547537
rect 0 546981 17809 546991
rect 0 546449 5481 546459
rect 0 545903 577836 546449
rect 0 545893 23053 545903
rect 0 545361 4101 545371
rect 0 544815 577836 545361
rect 0 544805 20753 544815
rect 0 544273 8793 544283
rect 0 543727 577836 544273
rect 0 543717 30781 543727
rect 0 543185 42649 543195
rect 0 542639 577836 543185
rect 0 542629 81105 542639
rect 0 542097 11277 542107
rect 0 541551 577836 542097
rect 0 541541 32621 541551
rect 0 541009 5205 541019
rect 0 540463 577836 541009
rect 0 540453 18637 540463
rect 0 539921 7413 539931
rect 0 539375 577836 539921
rect 0 539365 35381 539375
rect 0 538833 1801 538843
rect 0 538287 577836 538833
rect 0 538277 22869 538287
rect 0 537745 5573 537755
rect 0 537199 577836 537745
rect 0 537189 15233 537199
rect 0 536657 94445 536667
rect 0 536111 577836 536657
rect 0 536101 78897 536111
rect 0 535569 65281 535579
rect 0 535023 577836 535569
rect 0 535013 138421 535023
rect 0 534481 62705 534491
rect 0 533935 577836 534481
rect 0 533925 71905 533935
rect 0 533393 39153 533403
rect 0 532847 577836 533393
rect 0 532837 18913 532847
rect 0 532305 5389 532315
rect 0 531759 577836 532305
rect 0 531749 31057 531759
rect 0 531217 9161 531227
rect 0 530671 577836 531217
rect 0 530661 25813 530671
rect 0 530129 5297 530139
rect 0 529583 577836 530129
rect 0 529573 19189 529583
rect 0 529041 5297 529051
rect 0 528495 577836 529041
rect 0 528485 25537 528495
rect 0 527953 7413 527963
rect 0 527407 577836 527953
rect 0 527397 11553 527407
rect 0 526865 4745 526875
rect 0 526319 577836 526865
rect 0 526309 23697 526319
rect 0 525777 43753 525787
rect 0 525231 577836 525777
rect 0 525221 17349 525231
rect 0 524689 4653 524699
rect 0 524143 577836 524689
rect 0 524133 25537 524143
rect 0 523601 13025 523611
rect 0 523055 577836 523601
rect 0 523045 53965 523055
rect 0 522513 7321 522523
rect 0 521967 577836 522513
rect 0 521957 4561 521967
rect 0 521425 5205 521435
rect 0 520879 577836 521425
rect 0 520869 58105 520879
rect 0 520337 93433 520347
rect 0 519791 577836 520337
rect 0 519781 39613 519791
rect 0 519249 11369 519259
rect 0 518703 577836 519249
rect 0 518693 8517 518703
rect 0 518161 26365 518171
rect 0 517615 577836 518161
rect 0 517605 5941 517615
rect 0 517073 5665 517083
rect 0 516527 577836 517073
rect 0 516517 23973 516527
rect 0 515985 46145 515995
rect 0 515439 577836 515985
rect 0 515429 83129 515439
rect 0 514897 5297 514907
rect 0 514351 577836 514897
rect 0 514341 88557 514351
rect 0 513809 21581 513819
rect 0 513263 577836 513809
rect 0 513253 4561 513263
rect 0 512721 28297 512731
rect 0 512175 577836 512721
rect 0 512165 13393 512175
rect 0 511633 5113 511643
rect 0 511087 577836 511633
rect 0 511077 8701 511087
rect 0 510545 78621 510555
rect 0 509999 577836 510545
rect 0 509989 7689 509999
rect 0 509457 11277 509467
rect 0 508911 577836 509457
rect 0 508901 35013 508911
rect 0 508369 4929 508379
rect 0 507823 577836 508369
rect 0 507813 43845 507823
rect 0 507281 27285 507291
rect 0 506735 577836 507281
rect 0 506725 11553 506735
rect 0 506193 4653 506203
rect 0 505647 577836 506193
rect 0 505637 60589 505647
rect 0 505105 57645 505115
rect 0 504559 577836 505105
rect 0 504549 4561 504559
rect 0 504017 17533 504027
rect 0 503471 577836 504017
rect 0 503461 10173 503471
rect 0 502929 21029 502939
rect 0 502383 577836 502929
rect 0 502373 4561 502383
rect 0 501841 35473 501851
rect 0 501295 577836 501841
rect 0 501285 86993 501295
rect 0 500753 130509 500763
rect 0 500207 577836 500753
rect 0 500197 115053 500207
rect 0 499665 265013 499675
rect 0 499119 577836 499665
rect 0 499109 10173 499119
rect 0 498577 53781 498587
rect 0 498031 577836 498577
rect 0 498021 15785 498031
rect 0 497489 881 497499
rect 0 496943 577836 497489
rect 0 496933 3825 496943
rect 0 496401 23513 496411
rect 0 495855 577836 496401
rect 0 495845 14221 495855
rect 0 495313 59301 495323
rect 0 494767 577836 495313
rect 0 494757 4101 494767
rect 0 494225 16889 494235
rect 0 493679 577836 494225
rect 0 493669 52309 493679
rect 0 493137 881 493147
rect 0 492591 577836 493137
rect 0 492581 7597 492591
rect 0 492049 44857 492059
rect 0 491503 577836 492049
rect 0 491493 4561 491503
rect 0 490961 36853 490971
rect 0 490415 577836 490961
rect 0 490405 697 490415
rect 0 489873 28205 489883
rect 0 489327 577836 489873
rect 0 489317 7505 489327
rect 0 488785 4285 488795
rect 0 488239 577836 488785
rect 0 488229 789 488239
rect 0 487697 17625 487707
rect 0 487151 577836 487697
rect 0 487141 13945 487151
rect 0 486609 26089 486619
rect 0 486063 577836 486609
rect 0 486053 32161 486063
rect 0 485521 8977 485531
rect 0 484975 577836 485521
rect 0 484965 42189 484975
rect 0 484433 789 484443
rect 0 483887 577836 484433
rect 0 483877 4561 483887
rect 0 483345 24249 483355
rect 0 482799 577836 483345
rect 0 482789 68317 482799
rect 0 482257 18545 482267
rect 0 481711 577836 482257
rect 0 481701 31241 481711
rect 0 481169 84141 481179
rect 0 480623 577836 481169
rect 0 480613 3733 480623
rect 0 480081 1065 480091
rect 0 479535 577836 480081
rect 0 479525 24249 479535
rect 0 478993 15141 479003
rect 0 478447 577836 478993
rect 0 478437 81381 478447
rect 0 477905 12381 477915
rect 0 477359 577836 477905
rect 0 477349 4561 477359
rect 0 476817 24157 476827
rect 0 476271 577836 476817
rect 0 476261 8425 476271
rect 0 475729 1249 475739
rect 0 475183 577836 475729
rect 0 475173 112569 475183
rect 0 474641 12289 474651
rect 0 474095 577836 474641
rect 0 474085 43293 474095
rect 0 473553 8885 473563
rect 0 473007 577836 473553
rect 0 472997 2077 473007
rect 0 472465 5389 472475
rect 0 471919 577836 472465
rect 0 471909 53505 471919
rect 0 471377 17901 471387
rect 0 470831 577836 471377
rect 0 470821 37773 470831
rect 0 470289 4653 470299
rect 0 469743 577836 470289
rect 0 469733 8149 469743
rect 0 469201 24249 469211
rect 0 468655 577836 469201
rect 0 468645 697 468655
rect 0 468113 18637 468123
rect 0 467567 577836 468113
rect 0 467557 28481 467567
rect 0 467025 91501 467035
rect 0 466479 577836 467025
rect 0 466469 32345 466479
rect 0 465937 35105 465947
rect 0 465391 577836 465937
rect 0 465381 15785 465391
rect 0 464849 789 464859
rect 0 464303 577836 464849
rect 0 464293 3825 464303
rect 0 463761 10633 463771
rect 0 463215 577836 463761
rect 0 463205 7597 463215
rect 0 462673 1709 462683
rect 0 462127 577836 462673
rect 0 462117 67673 462127
rect 0 461585 100241 461595
rect 0 461039 577836 461585
rect 0 461029 88741 461039
rect 0 460497 61049 460507
rect 0 459951 577836 460497
rect 0 459941 135017 459951
rect 0 459409 16981 459419
rect 0 458863 577836 459409
rect 0 458853 513 458863
rect 0 458321 14405 458331
rect 0 457775 577836 458321
rect 0 457765 8609 457775
rect 0 457233 5573 457243
rect 0 456687 577836 457233
rect 0 456677 8793 456687
rect 0 456145 29861 456155
rect 0 455599 577836 456145
rect 0 455589 26641 455599
rect 0 455057 3181 455067
rect 0 454511 577836 455057
rect 0 454501 23329 454511
rect 0 453969 5757 453979
rect 0 453423 577836 453969
rect 0 453413 29953 453423
rect 0 452881 14865 452891
rect 0 452335 577836 452881
rect 0 452325 2169 452335
rect 0 451793 9621 451803
rect 0 451247 577836 451793
rect 0 451237 27009 451247
rect 0 450705 14405 450715
rect 0 450159 577836 450705
rect 0 450149 17257 450159
rect 0 449617 57921 449627
rect 0 449071 577836 449617
rect 0 449061 1157 449071
rect 0 448529 7413 448539
rect 0 447983 577836 448529
rect 0 447973 4469 447983
rect 0 447441 66385 447451
rect 0 446895 577836 447441
rect 0 446885 17441 446895
rect 0 446353 1341 446363
rect 0 445807 577836 446353
rect 0 445797 66293 445807
rect 0 445265 14497 445275
rect 0 444719 577836 445265
rect 0 444709 7965 444719
rect 0 444177 5113 444187
rect 0 443631 577836 444177
rect 0 443621 26641 443631
rect 0 443089 20201 443099
rect 0 442543 577836 443089
rect 0 442533 69145 442543
rect 0 442001 52217 442011
rect 0 441455 577836 442001
rect 0 441445 789 441455
rect 0 440913 29585 440923
rect 0 440367 577836 440913
rect 0 440357 68041 440367
rect 0 439825 10817 439835
rect 0 439279 577836 439825
rect 0 439269 1709 439279
rect 0 438737 42925 438747
rect 0 438191 577836 438737
rect 0 438181 4561 438191
rect 0 437649 13025 437659
rect 0 437103 577836 437649
rect 0 437093 26733 437103
rect 0 436561 55253 436571
rect 0 436015 577836 436561
rect 0 436005 9897 436015
rect 0 435473 18637 435483
rect 0 434927 577836 435473
rect 0 434917 973 434927
rect 0 434385 32989 434395
rect 0 433839 577836 434385
rect 0 433829 23053 433839
rect 0 433297 15049 433307
rect 0 432751 577836 433297
rect 0 432741 4561 432751
rect 0 432209 1801 432219
rect 0 431663 577836 432209
rect 0 431653 48353 431663
rect 0 431121 32989 431131
rect 0 430575 577836 431121
rect 0 430565 28941 430575
rect 0 430033 8793 430043
rect 0 429487 577836 430033
rect 0 429477 24617 429487
rect 0 428945 11553 428955
rect 0 428399 577836 428945
rect 0 428389 4285 428399
rect 0 427857 1801 427867
rect 0 427311 577836 427857
rect 0 427301 7413 427311
rect 0 426769 122597 426779
rect 0 426223 577836 426769
rect 0 426213 47617 426223
rect 0 425681 46697 425691
rect 0 425135 577836 425681
rect 0 425125 75217 425135
rect 0 424593 63073 424603
rect 0 424047 577836 424593
rect 0 424037 55069 424047
rect 0 423505 49917 423515
rect 0 422959 577836 423505
rect 0 422949 19373 422959
rect 0 422417 33357 422427
rect 0 421871 577836 422417
rect 0 421861 15785 421871
rect 0 421329 22501 421339
rect 0 420783 577836 421329
rect 0 420773 25537 420783
rect 0 420241 28941 420251
rect 0 419695 577836 420241
rect 0 419685 6585 419695
rect 0 419153 9897 419163
rect 0 418607 577836 419153
rect 0 418597 46697 418607
rect 0 418065 55621 418075
rect 0 417519 577836 418065
rect 0 417509 1065 417519
rect 0 416977 8977 416987
rect 0 416431 577836 416977
rect 0 416421 34001 416431
rect 0 415889 12381 415899
rect 0 415343 577836 415889
rect 0 415333 19557 415343
rect 0 414801 67673 414811
rect 0 414255 577836 414801
rect 0 414245 82761 414255
rect 0 413713 16153 413723
rect 0 413167 577836 413713
rect 0 413157 881 413167
rect 0 412625 5941 412635
rect 0 412079 577836 412625
rect 0 412069 25077 412079
rect 0 411537 9897 411547
rect 0 410991 577836 411537
rect 0 410981 12565 410991
rect 0 410449 72733 410459
rect 0 409903 577836 410449
rect 0 409893 92513 409903
rect 0 409361 3733 409371
rect 0 408815 577836 409361
rect 0 408805 1341 408815
rect 0 408273 18269 408283
rect 0 407727 577836 408273
rect 0 407717 30781 407727
rect 0 407185 27745 407195
rect 0 406639 577836 407185
rect 0 406629 41361 406639
rect 0 406097 24249 406107
rect 0 405551 577836 406097
rect 0 405541 973 405551
rect 0 405009 21581 405019
rect 0 404463 577836 405009
rect 0 404453 19097 404463
rect 0 403921 50837 403931
rect 0 403375 577836 403921
rect 0 403365 2721 403375
rect 0 402833 27561 402843
rect 0 402287 577836 402833
rect 0 402277 6493 402287
rect 0 401745 31517 401755
rect 0 401199 577836 401745
rect 0 401189 789 401199
rect 0 400657 21857 400667
rect 0 400111 577836 400657
rect 0 400101 5941 400111
rect 0 399569 7229 399579
rect 0 399023 577836 399569
rect 0 399013 10173 399023
rect 0 398481 18637 398491
rect 0 397935 577836 398481
rect 0 397925 2537 397935
rect 0 397393 9621 397403
rect 0 396847 577836 397393
rect 0 396837 1985 396847
rect 0 396305 3181 396315
rect 0 395759 577836 396305
rect 0 395749 6493 395759
rect 0 395217 29861 395227
rect 0 394671 577836 395217
rect 0 394661 167309 394671
rect 0 394129 13025 394139
rect 0 393583 577836 394129
rect 0 393573 1249 393583
rect 0 393041 17901 393051
rect 0 392495 577836 393041
rect 0 392485 4377 392495
rect 0 391953 37405 391963
rect 0 391407 577836 391953
rect 0 391397 7505 391407
rect 0 390865 34645 390875
rect 0 390319 577836 390865
rect 0 390309 10173 390319
rect 0 389777 1341 389787
rect 0 389231 577836 389777
rect 0 389221 14221 389231
rect 0 388689 4469 388699
rect 0 388143 577836 388689
rect 0 388133 7965 388143
rect 0 387601 37221 387611
rect 0 387055 577836 387601
rect 0 387045 18729 387055
rect 0 386513 74757 386523
rect 0 385967 577836 386513
rect 0 385957 13025 385967
rect 0 385425 1249 385435
rect 0 384879 577836 385425
rect 0 384869 38233 384879
rect 0 384337 28021 384347
rect 0 383791 577836 384337
rect 0 383781 2537 383791
rect 0 383249 18637 383259
rect 0 382703 577836 383249
rect 0 382693 63717 382703
rect 0 382161 13025 382171
rect 0 381615 577836 382161
rect 0 381605 10081 381615
rect 0 381073 74389 381083
rect 0 380527 577836 381073
rect 0 380517 49089 380527
rect 0 379985 8793 379995
rect 0 379439 577836 379985
rect 0 379429 24433 379439
rect 0 378897 12933 378907
rect 0 378351 577836 378897
rect 0 378341 2169 378351
rect 0 377809 21029 377819
rect 0 377263 577836 377809
rect 0 377253 41545 377263
rect 0 376721 9345 376731
rect 0 376175 577836 376721
rect 0 376165 3549 376175
rect 0 375633 4929 375643
rect 0 375087 577836 375633
rect 0 375077 30689 375087
rect 0 374545 48261 374555
rect 0 373999 577836 374545
rect 0 373989 18913 373999
rect 0 373457 6033 373467
rect 0 372911 577836 373457
rect 0 372901 7413 372911
rect 0 372369 10725 372379
rect 0 371823 577836 372369
rect 0 371813 69605 371823
rect 0 371281 32805 371291
rect 0 370735 577836 371281
rect 0 370725 35749 370735
rect 0 370193 18637 370203
rect 0 369647 577836 370193
rect 0 369637 3089 369647
rect 0 369105 3181 369115
rect 0 368559 577836 369105
rect 0 368549 7965 368559
rect 0 368017 15509 368027
rect 0 367471 577836 368017
rect 0 367461 4561 367471
rect 0 366929 3917 366939
rect 0 366383 577836 366929
rect 0 366373 35473 366383
rect 0 365841 7413 365851
rect 0 365295 577836 365841
rect 0 365285 32161 365295
rect 0 364753 3181 364763
rect 0 364207 577836 364753
rect 0 364197 17165 364207
rect 0 363665 26733 363675
rect 0 363119 577836 363665
rect 0 363109 110913 363119
rect 0 362577 4469 362587
rect 0 362031 577836 362577
rect 0 362021 3089 362031
rect 0 361489 16337 361499
rect 0 360943 577836 361489
rect 0 360933 32621 360943
rect 0 360401 28205 360411
rect 0 359855 577836 360401
rect 0 359845 76873 359855
rect 0 359313 1525 359323
rect 0 358767 577836 359313
rect 0 358757 65649 358767
rect 0 358225 4653 358235
rect 0 357679 577836 358225
rect 0 357669 10173 357679
rect 0 357137 7413 357147
rect 0 356591 577836 357137
rect 0 356581 34093 356591
rect 0 356049 22225 356059
rect 0 355503 577836 356049
rect 0 355493 76965 355503
rect 0 354961 85981 354971
rect 0 354415 577836 354961
rect 0 354405 66293 354415
rect 0 353873 105761 353883
rect 0 353327 577836 353873
rect 0 353317 60681 353327
rect 0 352785 107877 352795
rect 0 352239 577836 352785
rect 0 352229 63533 352239
rect 0 351697 67673 351707
rect 0 351151 577836 351697
rect 0 351141 4285 351151
rect 0 350609 209261 350619
rect 0 350063 577836 350609
rect 0 350053 23053 350063
rect 0 349521 3181 349531
rect 0 348975 577836 349521
rect 0 348965 11829 348975
rect 0 348433 8793 348443
rect 0 347887 577836 348433
rect 0 347877 36209 347887
rect 0 347345 34369 347355
rect 0 346799 577836 347345
rect 0 346789 43569 346799
rect 0 346257 33725 346267
rect 0 345711 577836 346257
rect 0 345701 4285 345711
rect 0 345169 3181 345179
rect 0 344623 577836 345169
rect 0 344613 32621 344623
rect 0 344081 12933 344091
rect 0 343535 577836 344081
rect 0 343525 38049 343535
rect 0 342993 9897 343003
rect 0 342447 577836 342993
rect 0 342437 6861 342447
rect 0 341905 12473 341915
rect 0 341359 577836 341905
rect 0 341349 3917 341359
rect 0 340817 18361 340827
rect 0 340271 577836 340817
rect 0 340261 29953 340271
rect 0 339729 27745 339739
rect 0 339183 577836 339729
rect 0 339173 85153 339183
rect 0 338641 3365 338651
rect 0 338095 577836 338641
rect 0 338085 21397 338095
rect 0 337553 12013 337563
rect 0 337007 577836 337553
rect 0 336997 15785 337007
rect 0 336465 8793 336475
rect 0 335919 577836 336465
rect 0 335909 64637 335919
rect 0 335377 11553 335387
rect 0 334831 577836 335377
rect 0 334821 36669 334831
rect 0 334289 3365 334299
rect 0 333743 577836 334289
rect 0 333733 28849 333743
rect 0 333201 42833 333211
rect 0 332655 577836 333201
rect 0 332645 8333 332655
rect 0 332113 14405 332123
rect 0 331567 577836 332113
rect 0 331557 23145 331567
rect 0 331025 3457 331035
rect 0 330479 577836 331025
rect 0 330469 42465 330479
rect 0 329937 64913 329947
rect 0 329391 577836 329937
rect 0 329381 7597 329391
rect 0 328849 45133 328859
rect 0 328303 577836 328849
rect 0 328293 22777 328303
rect 0 327761 5389 327771
rect 0 327215 577836 327761
rect 0 327205 3365 327215
rect 0 326673 10265 326683
rect 0 326127 577836 326673
rect 0 326117 4193 326127
rect 0 325585 6309 325595
rect 0 325039 577836 325585
rect 0 325029 17717 325039
rect 0 324497 385257 324507
rect 0 323951 577836 324497
rect 0 323941 38233 323951
rect 0 323409 25905 323419
rect 0 322863 577836 323409
rect 0 322853 4193 322863
rect 0 322321 9529 322331
rect 0 321775 577836 322321
rect 0 321765 47893 321775
rect 0 321233 7137 321243
rect 0 320687 577836 321233
rect 0 320677 4193 320687
rect 0 320145 18545 320155
rect 0 319599 577836 320145
rect 0 319589 23237 319599
rect 0 319057 97205 319067
rect 0 318511 577836 319057
rect 0 318501 28389 318511
rect 0 317969 6769 317979
rect 0 317423 577836 317969
rect 0 317413 3825 317423
rect 0 316881 34461 316891
rect 0 316335 577836 316881
rect 0 316325 9897 316335
rect 0 315793 15141 315803
rect 0 315247 577836 315793
rect 0 315237 31149 315247
rect 0 314705 28941 314715
rect 0 314159 577836 314705
rect 0 314149 60037 314159
rect 0 313617 4653 313627
rect 0 313071 577836 313617
rect 0 313061 22777 313071
rect 0 312529 12657 312539
rect 0 311983 577836 312529
rect 0 311973 29953 311983
rect 0 311441 15417 311451
rect 0 310895 577836 311441
rect 0 310885 4193 310895
rect 0 310353 12013 310363
rect 0 309807 577836 310353
rect 0 309797 32069 309807
rect 0 309265 24157 309275
rect 0 308719 577836 309265
rect 0 308709 71905 308719
rect 0 308177 82393 308187
rect 0 307631 577836 308177
rect 0 307621 18913 307631
rect 0 307089 6585 307099
rect 0 306543 577836 307089
rect 0 306533 3457 306543
rect 0 306001 15877 306011
rect 0 305455 577836 306001
rect 0 305445 31149 305455
rect 0 304913 31241 304923
rect 0 304367 577836 304913
rect 0 304357 4101 304367
rect 0 303825 6677 303835
rect 0 303279 577836 303825
rect 0 303269 13025 303279
rect 0 302737 21673 302747
rect 0 302191 577836 302737
rect 0 302181 84509 302191
rect 0 301649 15877 301659
rect 0 301103 577836 301649
rect 0 301093 24525 301103
rect 0 300561 10265 300571
rect 0 300015 577836 300561
rect 0 300005 90121 300015
rect 0 299473 13025 299483
rect 0 298927 577836 299473
rect 0 298917 6493 298927
rect 0 298385 10081 298395
rect 0 297839 577836 298385
rect 0 297829 32621 297839
rect 0 297297 5297 297307
rect 0 296751 577836 297297
rect 0 296741 19097 296751
rect 0 296209 14405 296219
rect 0 295663 577836 296209
rect 0 295653 34001 295663
rect 0 295121 9529 295131
rect 0 294575 577836 295121
rect 0 294565 4009 294575
rect 0 294033 22225 294043
rect 0 293487 577836 294033
rect 0 293477 36669 293487
rect 0 292945 66753 292955
rect 0 292399 577836 292945
rect 0 292389 17809 292399
rect 0 291857 13025 291867
rect 0 291311 577836 291857
rect 0 291301 23421 291311
rect 0 290769 11461 290779
rect 0 290223 577836 290769
rect 0 290213 19557 290223
rect 0 289681 114041 289691
rect 0 289135 577836 289681
rect 0 289125 65005 289135
rect 0 288593 66661 288603
rect 0 288047 577836 288593
rect 0 288037 75861 288047
rect 0 287505 73285 287515
rect 0 286959 577836 287505
rect 0 286949 70617 286959
rect 0 286417 48261 286427
rect 0 285871 577836 286417
rect 0 285861 25077 285871
rect 0 285329 9345 285339
rect 0 284783 577836 285329
rect 0 284773 15785 284783
rect 0 284241 21765 284251
rect 0 283695 577836 284241
rect 0 283685 28757 283695
rect 0 283153 39613 283163
rect 0 282607 577836 283153
rect 0 282597 12473 282607
rect 0 282065 98861 282075
rect 0 281519 577836 282065
rect 0 281509 41637 281519
rect 0 280977 12565 280987
rect 0 280431 577836 280977
rect 0 280421 6125 280431
rect 0 279889 6033 279899
rect 0 279343 577836 279889
rect 0 279333 9989 279343
rect 0 278801 49549 278811
rect 0 278255 577836 278801
rect 0 278245 15049 278255
rect 0 277713 29769 277723
rect 0 277167 577836 277713
rect 0 277157 11645 277167
rect 0 276625 3917 276635
rect 0 276079 577836 276625
rect 0 276069 17717 276079
rect 0 275537 24249 275547
rect 0 274991 577836 275537
rect 0 274981 4009 274991
rect 0 274449 18637 274459
rect 0 273903 577836 274449
rect 0 273893 8609 273903
rect 0 273361 33541 273371
rect 0 272815 577836 273361
rect 0 272805 2445 272815
rect 0 272273 11553 272283
rect 0 271727 577836 272273
rect 0 271717 14957 271727
rect 0 271185 12013 271195
rect 0 270639 577836 271185
rect 0 270629 42281 270639
rect 0 270097 39061 270107
rect 0 269551 577836 270097
rect 0 269541 2813 269551
rect 0 269009 29861 269019
rect 0 268463 577836 269009
rect 0 268453 9069 268463
rect 0 267921 18637 267931
rect 0 267375 577836 267921
rect 0 267365 57829 267375
rect 0 266833 139341 266843
rect 0 266287 577836 266833
rect 0 266277 2905 266287
rect 0 265745 70525 265755
rect 0 265199 577836 265745
rect 0 265189 21397 265199
rect 0 264657 9713 264667
rect 0 264111 577836 264657
rect 0 264101 54701 264111
rect 0 263569 17717 263579
rect 0 263023 577836 263569
rect 0 263013 5941 263023
rect 0 262481 69145 262491
rect 0 261935 577836 262481
rect 0 261925 5941 261935
rect 0 261393 124621 261403
rect 0 260847 577836 261393
rect 0 260837 103645 260847
rect 0 260305 18545 260315
rect 0 259759 577836 260305
rect 0 259749 15785 259759
rect 0 259217 26089 259227
rect 0 258671 577836 259217
rect 0 258661 5941 258671
rect 0 258129 12105 258139
rect 0 257583 577836 258129
rect 0 257573 3917 257583
rect 0 257041 12473 257051
rect 0 256495 577836 257041
rect 0 256485 40073 256495
rect 0 255953 29309 255963
rect 0 255407 577836 255953
rect 0 255397 8977 255407
rect 0 254865 14405 254875
rect 0 254319 577836 254865
rect 0 254309 15693 254319
rect 0 253777 5297 253787
rect 0 253231 577836 253777
rect 0 253221 8149 253231
rect 0 252689 42465 252699
rect 0 252143 577836 252689
rect 0 252133 13393 252143
rect 0 251601 23697 251611
rect 0 251055 577836 251601
rect 0 251045 17165 251055
rect 0 250513 49549 250523
rect 0 249967 577836 250513
rect 0 249957 2537 249967
rect 0 249425 5573 249435
rect 0 248879 577836 249425
rect 0 248869 40349 248879
rect 0 248337 59301 248347
rect 0 247791 577836 248337
rect 0 247781 15785 247791
rect 0 247249 43937 247259
rect 0 246703 577836 247249
rect 0 246693 18913 246703
rect 0 246161 10541 246171
rect 0 245615 577836 246161
rect 0 245605 15049 245615
rect 0 245073 3825 245083
rect 0 244527 577836 245073
rect 0 244517 32345 244527
rect 0 243985 16061 243995
rect 0 243439 577836 243985
rect 0 243429 4561 243439
rect 0 242897 48169 242907
rect 0 242351 577836 242897
rect 0 242341 27009 242351
rect 0 241809 10541 241819
rect 0 241263 577836 241809
rect 0 241253 14865 241263
rect 0 240721 6769 240731
rect 0 240175 577836 240721
rect 0 240165 18729 240175
rect 0 239633 24249 239643
rect 0 239087 577836 239633
rect 0 239077 3181 239087
rect 0 238545 27653 238555
rect 0 237999 577836 238545
rect 0 237989 13301 237999
rect 0 237457 9345 237467
rect 0 236911 577836 237457
rect 0 236901 2905 236911
rect 0 236369 28389 236379
rect 0 235823 577836 236369
rect 0 235813 69513 235823
rect 0 235281 39797 235291
rect 0 234735 577836 235281
rect 0 234725 39613 234735
rect 0 234193 14405 234203
rect 0 233647 577836 234193
rect 0 233637 51941 233647
rect 0 233105 48629 233115
rect 0 232559 577836 233105
rect 0 232549 4469 232559
rect 0 232017 11185 232027
rect 0 231471 577836 232017
rect 0 231461 51665 231471
rect 0 230929 22133 230939
rect 0 230383 577836 230929
rect 0 230373 96009 230383
rect 0 229841 85981 229851
rect 0 229295 577836 229841
rect 0 229285 84969 229295
rect 0 228753 76137 228763
rect 0 228207 577836 228753
rect 0 228197 67857 228207
rect 0 227665 16521 227675
rect 0 227119 577836 227665
rect 0 227109 35105 227119
rect 0 226577 22685 226587
rect 0 226031 577836 226577
rect 0 226021 7597 226031
rect 0 225489 1617 225499
rect 0 224943 577836 225489
rect 0 224933 4469 224943
rect 0 224401 137869 224411
rect 0 223855 577836 224401
rect 0 223845 10173 223855
rect 0 223313 29861 223323
rect 0 222767 577836 223313
rect 0 222757 4469 222767
rect 0 222225 20017 222235
rect 0 221679 577836 222225
rect 0 221669 35749 221679
rect 0 221137 10541 221147
rect 0 220591 577836 221137
rect 0 220581 2077 220591
rect 0 220049 4193 220059
rect 0 219503 577836 220049
rect 0 219493 26825 219503
rect 0 218961 1801 218971
rect 0 218415 577836 218961
rect 0 218405 71077 218415
rect 0 217873 15417 217883
rect 0 217327 577836 217873
rect 0 217317 9345 217327
rect 0 216785 29861 216795
rect 0 216239 577836 216785
rect 0 216229 43017 216239
rect 0 215697 1801 215707
rect 0 215151 577836 215697
rect 0 215141 41085 215151
rect 0 214609 11277 214619
rect 0 214063 577836 214609
rect 0 214053 15601 214063
rect 0 213521 5941 213531
rect 0 212975 577836 213521
rect 0 212965 77517 212975
rect 0 212433 8793 212443
rect 0 211887 577836 212433
rect 0 211877 28389 211887
rect 0 211345 16429 211355
rect 0 210799 577836 211345
rect 0 210789 10173 210799
rect 0 210257 7413 210267
rect 0 209711 577836 210257
rect 0 209701 1249 209711
rect 0 209169 29401 209179
rect 0 208623 577836 209169
rect 0 208613 15417 208623
rect 0 208081 5389 208091
rect 0 207535 577836 208081
rect 0 207525 13117 207535
rect 0 206993 1433 207003
rect 0 206447 577836 206993
rect 0 206437 22777 206447
rect 0 205905 15417 205915
rect 0 205359 577836 205905
rect 0 205349 108613 205359
rect 0 204817 29125 204827
rect 0 204271 577836 204817
rect 0 204261 13853 204271
rect 0 203729 1617 203739
rect 0 203183 577836 203729
rect 0 203173 9345 203183
rect 0 202641 4745 202651
rect 0 202095 577836 202641
rect 0 202085 36669 202095
rect 0 201553 1801 201563
rect 0 201007 577836 201553
rect 0 200997 30597 201007
rect 0 200465 40901 200475
rect 0 199919 577836 200465
rect 0 199909 14129 199919
rect 0 199377 11093 199387
rect 0 198831 577836 199377
rect 0 198821 7873 198831
rect 0 198289 4745 198299
rect 0 197743 577836 198289
rect 0 197733 46973 197743
rect 0 197201 39429 197211
rect 0 196655 577836 197201
rect 0 196645 83037 196655
rect 0 196113 1525 196123
rect 0 195567 577836 196113
rect 0 195557 13945 195567
rect 0 195025 42465 195035
rect 0 194479 577836 195025
rect 0 194469 8149 194479
rect 0 193937 1709 193947
rect 0 193391 577836 193937
rect 0 193381 17165 193391
rect 0 192849 36853 192859
rect 0 192303 577836 192849
rect 0 192293 1341 192303
rect 0 191761 17165 191771
rect 0 191215 577836 191761
rect 0 191205 43845 191215
rect 0 190673 11645 190683
rect 0 190127 577836 190673
rect 0 190117 4561 190127
rect 0 189585 48353 189595
rect 0 189039 577836 189585
rect 0 189029 103093 189039
rect 0 188497 3457 188507
rect 0 187951 577836 188497
rect 0 187941 17349 187951
rect 0 187409 11093 187419
rect 0 186863 577836 187409
rect 0 186853 74021 186863
rect 0 186321 1801 186331
rect 0 185775 577836 186321
rect 0 185765 7781 185775
rect 0 185233 33633 185243
rect 0 184687 577836 185233
rect 0 184677 77425 184687
rect 0 184145 10449 184155
rect 0 183599 577836 184145
rect 0 183589 15785 183599
rect 0 183057 3273 183067
rect 0 182511 577836 183057
rect 0 182501 24617 182511
rect 0 181969 74665 181979
rect 0 181423 577836 181969
rect 0 181413 10173 181423
rect 0 180881 20937 180891
rect 0 180335 577836 180881
rect 0 180325 1617 180335
rect 0 179793 6861 179803
rect 0 179247 577836 179793
rect 0 179237 46697 179247
rect 0 178705 16337 178715
rect 0 178159 577836 178705
rect 0 178149 38233 178159
rect 0 177617 13025 177627
rect 0 177071 577836 177617
rect 0 177061 9713 177071
rect 0 176529 3641 176539
rect 0 175983 577836 176529
rect 0 175973 17165 175983
rect 0 175441 20201 175451
rect 0 174895 577836 175441
rect 0 174885 29677 174895
rect 0 174353 40717 174363
rect 0 173807 577836 174353
rect 0 173797 88373 173807
rect 0 173265 13025 173275
rect 0 172719 577836 173265
rect 0 172709 64821 172719
rect 0 172177 31241 172187
rect 0 171631 577836 172177
rect 0 171621 22869 171631
rect 0 171089 16797 171099
rect 0 170543 577836 171089
rect 0 170533 43109 170543
rect 0 170001 42833 170011
rect 0 169455 577836 170001
rect 0 169445 88741 169455
rect 0 168913 39429 168923
rect 0 168367 577836 168913
rect 0 168357 50837 168367
rect 0 167825 60773 167835
rect 0 167279 577836 167825
rect 0 167269 26825 167279
rect 0 166737 14497 166747
rect 0 166191 577836 166737
rect 0 166181 2813 166191
rect 0 165649 513 165659
rect 0 165103 577836 165649
rect 0 165093 5941 165103
rect 0 164561 27929 164571
rect 0 164015 577836 164561
rect 0 164005 12013 164015
rect 0 163473 7045 163483
rect 0 162927 577836 163473
rect 0 162917 36761 162927
rect 0 162385 63257 162395
rect 0 161839 577836 162385
rect 0 161829 9897 161839
rect 0 161297 42649 161307
rect 0 160751 577836 161297
rect 0 160741 15509 160751
rect 0 160209 1709 160219
rect 0 159663 577836 160209
rect 0 159653 4469 159663
rect 0 159121 126829 159131
rect 0 158575 577836 159121
rect 0 158565 35749 158575
rect 0 158033 32989 158043
rect 0 157487 577836 158033
rect 0 157477 12289 157487
rect 0 156945 17901 156955
rect 0 156399 577836 156945
rect 0 156389 22961 156399
rect 0 155857 8793 155867
rect 0 155311 577836 155857
rect 0 155301 8517 155311
rect 0 154769 1801 154779
rect 0 154223 577836 154769
rect 0 154213 11829 154223
rect 0 153681 36945 153691
rect 0 153135 577836 153681
rect 0 153125 15785 153135
rect 0 152593 51665 152603
rect 0 152047 577836 152593
rect 0 152037 3089 152047
rect 0 151505 605 151515
rect 0 150959 577836 151505
rect 0 150949 6585 150959
rect 0 150417 22133 150427
rect 0 149871 577836 150417
rect 0 149861 54517 149871
rect 0 149329 3181 149339
rect 0 148783 577836 149329
rect 0 148773 18913 148783
rect 0 148241 13025 148251
rect 0 147695 577836 148241
rect 0 147685 67673 147695
rect 0 147153 42649 147163
rect 0 146607 577836 147153
rect 0 146597 39981 146607
rect 0 146065 6217 146075
rect 0 145519 577836 146065
rect 0 145509 152221 145519
rect 0 144977 29769 144987
rect 0 144431 577836 144977
rect 0 144421 42741 144431
rect 0 143889 1525 143899
rect 0 143343 577836 143889
rect 0 143333 11553 143343
rect 0 142801 37865 142811
rect 0 142255 577836 142801
rect 0 142245 2813 142255
rect 0 141713 8793 141723
rect 0 141167 577836 141713
rect 0 141157 42097 141167
rect 0 140625 5573 140635
rect 0 140079 577836 140625
rect 0 140069 56449 140079
rect 0 139537 65833 139547
rect 0 138991 577836 139537
rect 0 138981 2445 138991
rect 0 138449 8793 138459
rect 0 137903 577836 138449
rect 0 137893 37037 137903
rect 0 137361 5113 137371
rect 0 136815 577836 137361
rect 0 136805 513 136815
rect 0 136273 17073 136283
rect 0 135727 577836 136273
rect 0 135717 14037 135727
rect 0 135185 56173 135195
rect 0 134639 577836 135185
rect 0 134629 8517 134639
rect 0 134097 513 134107
rect 0 133551 577836 134097
rect 0 133541 41913 133551
rect 0 133009 25629 133019
rect 0 132463 577836 133009
rect 0 132453 2997 132463
rect 0 131921 3181 131931
rect 0 131375 577836 131921
rect 0 131365 6217 131375
rect 0 130833 81749 130843
rect 0 130287 577836 130833
rect 0 130277 15233 130287
rect 0 129745 33173 129755
rect 0 129199 577836 129745
rect 0 129189 513 129199
rect 0 128657 11553 128667
rect 0 128111 577836 128657
rect 0 128101 14221 128111
rect 0 127569 46605 127579
rect 0 127023 577836 127569
rect 0 127013 32621 127023
rect 0 126481 20017 126491
rect 0 125935 577836 126481
rect 0 125925 36669 125935
rect 0 125393 93525 125403
rect 0 124847 577836 125393
rect 0 124837 11921 124847
rect 0 124305 7321 124315
rect 0 123759 577836 124305
rect 0 123749 513 123759
rect 0 123217 41085 123227
rect 0 122671 577836 123217
rect 0 122661 19465 122671
rect 0 122129 9161 122139
rect 0 121583 577836 122129
rect 0 121573 3825 121583
rect 0 121041 28205 121051
rect 0 120495 577836 121041
rect 0 120485 15049 120495
rect 0 119953 18545 119963
rect 0 119407 577836 119953
rect 0 119397 38233 119407
rect 0 118865 11553 118875
rect 0 118319 577836 118865
rect 0 118309 513 118319
rect 0 117777 6953 117787
rect 0 117231 577836 117777
rect 0 117221 2813 117231
rect 0 116689 53689 116699
rect 0 116143 577836 116689
rect 0 116133 66293 116143
rect 0 115601 3365 115611
rect 0 115055 577836 115601
rect 0 115045 37957 115055
rect 0 114513 11829 114523
rect 0 113967 577836 114513
rect 0 113957 3457 113967
rect 0 113425 513 113435
rect 0 112879 577836 113425
rect 0 112869 24617 112879
rect 0 112337 8885 112347
rect 0 111791 577836 112337
rect 0 111781 31149 111791
rect 0 111249 36853 111259
rect 0 110703 577836 111249
rect 0 110693 31517 110703
rect 0 110161 15325 110171
rect 0 109615 577836 110161
rect 0 109605 10173 109615
rect 0 109073 27377 109083
rect 0 108527 577836 109073
rect 0 108517 1341 108527
rect 0 107985 23053 107995
rect 0 107439 577836 107985
rect 0 107429 2077 107439
rect 0 106897 49917 106907
rect 0 106351 577836 106897
rect 0 106341 8149 106351
rect 0 105809 57553 105819
rect 0 105263 577836 105809
rect 0 105253 513 105263
rect 0 104721 5573 104731
rect 0 104175 577836 104721
rect 0 104165 79357 104175
rect 0 103633 12013 103643
rect 0 103087 577836 103633
rect 0 103077 2445 103087
rect 0 102545 10817 102555
rect 0 101999 577836 102545
rect 0 101989 15049 101999
rect 0 101457 7413 101467
rect 0 100911 577836 101457
rect 0 100901 56633 100911
rect 0 100369 37773 100379
rect 0 99823 577836 100369
rect 0 99813 513 99823
rect 0 99281 7229 99291
rect 0 98735 577836 99281
rect 0 98725 49089 98735
rect 0 98193 1801 98203
rect 0 97647 577836 98193
rect 0 97637 9805 97647
rect 0 97105 1525 97115
rect 0 96559 577836 97105
rect 0 96549 14313 96559
rect 0 96017 46513 96027
rect 0 95471 577836 96017
rect 0 95461 8885 95471
rect 0 94929 5297 94939
rect 0 94383 577836 94929
rect 0 94373 11737 94383
rect 0 93841 28389 93851
rect 0 93295 577836 93841
rect 0 93285 22777 93295
rect 0 92753 38601 92763
rect 0 92207 577836 92753
rect 0 92197 18729 92207
rect 0 91665 11461 91675
rect 0 91119 577836 91665
rect 0 91109 37037 91119
rect 0 90577 7137 90587
rect 0 90031 577836 90577
rect 0 90021 7413 90031
rect 0 89489 513 89499
rect 0 88943 577836 89489
rect 0 88933 70525 88943
rect 0 88401 17809 88411
rect 0 87855 577836 88401
rect 0 87845 3089 87855
rect 0 87313 38693 87323
rect 0 86767 577836 87313
rect 0 86757 22869 86767
rect 0 86225 95089 86235
rect 0 85679 577836 86225
rect 0 85669 24433 85679
rect 0 85137 16337 85147
rect 0 84591 577836 85137
rect 0 84581 9805 84591
rect 0 84049 24249 84059
rect 0 83503 577836 84049
rect 0 83493 513 83503
rect 0 82961 41085 82971
rect 0 82415 577836 82961
rect 0 82405 45777 82415
rect 0 81873 1157 81883
rect 0 81327 577836 81873
rect 0 81317 34001 81327
rect 0 80785 90489 80795
rect 0 80239 577836 80785
rect 0 80229 22777 80239
rect 0 79697 8885 79707
rect 0 79151 577836 79697
rect 0 79141 4561 79151
rect 0 78609 10449 78619
rect 0 78063 577836 78609
rect 0 78053 2169 78063
rect 0 77521 10633 77531
rect 0 76975 577836 77521
rect 0 76965 513 76975
rect 0 76433 11829 76443
rect 0 75887 577836 76433
rect 0 75877 30505 75887
rect 0 75345 27101 75355
rect 0 74799 577836 75345
rect 0 74789 96101 74799
rect 0 74257 1801 74267
rect 0 73711 577836 74257
rect 0 73701 1617 73711
rect 0 73169 22041 73179
rect 0 72623 577836 73169
rect 0 72613 14129 72623
rect 0 72081 76137 72091
rect 0 71535 577836 72081
rect 0 71525 62061 71535
rect 0 70993 71077 71003
rect 0 70447 577836 70993
rect 0 70437 13761 70447
rect 0 69905 35473 69915
rect 0 69359 577836 69905
rect 0 69349 81289 69359
rect 0 68817 40901 68827
rect 0 68271 577836 68817
rect 0 68261 23145 68271
rect 0 67729 20937 67739
rect 0 67183 577836 67729
rect 0 67173 17625 67183
rect 0 66641 39245 66651
rect 0 66095 577836 66641
rect 0 66085 99965 66095
rect 0 65553 27837 65563
rect 0 65007 577836 65553
rect 0 64997 8701 65007
rect 0 64465 8793 64475
rect 0 63919 577836 64465
rect 0 63909 22777 63919
rect 0 63377 10265 63387
rect 0 62831 577836 63377
rect 0 62821 36117 62831
rect 0 62289 63441 62299
rect 0 61743 577836 62289
rect 0 61733 34553 61743
rect 0 61201 27101 61211
rect 0 60655 577836 61201
rect 0 60645 30597 60655
rect 0 60113 20477 60123
rect 0 59567 577836 60113
rect 0 59557 9805 59567
rect 0 59025 40165 59035
rect 0 58479 577836 59025
rect 0 58469 12657 58479
rect 0 57937 6769 57947
rect 0 57391 577836 57937
rect 0 57381 24249 57391
rect 0 56849 74389 56859
rect 0 56303 577836 56849
rect 0 56293 51665 56303
rect 0 55761 14405 55771
rect 0 55215 577836 55761
rect 0 55205 8241 55215
rect 0 54673 31241 54683
rect 0 54127 577836 54673
rect 0 54117 7505 54127
rect 0 53585 40349 53595
rect 0 53039 577836 53585
rect 0 53029 15325 53039
rect 0 52497 74757 52507
rect 0 51951 577836 52497
rect 0 51941 53413 51951
rect 0 51409 20017 51419
rect 0 50863 577836 51409
rect 0 50853 22961 50863
rect 0 50321 10265 50331
rect 0 49775 577836 50321
rect 0 49765 15141 49775
rect 0 49233 33449 49243
rect 0 48687 577836 49233
rect 0 48677 26089 48687
rect 0 48145 7413 48155
rect 0 47599 577836 48145
rect 0 47589 56633 47599
rect 0 47057 18637 47067
rect 0 46511 577836 47057
rect 0 46501 11921 46511
rect 0 45969 22409 45979
rect 0 45423 577836 45969
rect 0 45413 12197 45423
rect 0 44881 9253 44891
rect 0 44335 577836 44881
rect 0 44325 36025 44335
rect 0 43793 22593 43803
rect 0 43247 577836 43793
rect 0 43237 7413 43247
rect 0 42705 196749 42715
rect 0 42159 577836 42705
rect 0 42149 13117 42159
rect 0 41617 20201 41627
rect 0 41071 577836 41617
rect 0 41061 17349 41071
rect 0 40529 18085 40539
rect 0 39983 577836 40529
rect 0 39973 7413 39983
rect 0 39441 10541 39451
rect 0 38895 577836 39441
rect 0 38885 20845 38895
rect 0 38353 10541 38363
rect 0 37807 577836 38353
rect 0 37797 47893 37807
rect 0 37265 15877 37275
rect 0 36719 577836 37265
rect 0 36709 67673 36719
rect 0 36177 12657 36187
rect 0 35631 577836 36177
rect 0 35621 63533 35631
rect 0 35089 22685 35099
rect 0 34543 577836 35089
rect 0 34533 50837 34543
rect 0 34001 35289 34011
rect 0 33455 577836 34001
rect 0 33445 39613 33455
rect 0 32913 20017 32923
rect 0 32367 577836 32913
rect 0 32357 31977 32367
rect 0 31825 17625 31835
rect 0 31279 577836 31825
rect 0 31269 7965 31279
rect 0 30737 39061 30747
rect 0 30191 577836 30737
rect 0 30181 50837 30191
rect 0 29649 43477 29659
rect 0 29103 577836 29649
rect 0 29093 26549 29103
rect 0 28561 34645 28571
rect 0 28015 577836 28561
rect 0 28005 17809 28015
rect 0 27473 61969 27483
rect 0 26927 577836 27473
rect 0 26917 9529 26927
rect 0 26385 18177 26395
rect 0 25839 577836 26385
rect 0 25829 17717 25839
rect 0 25297 224533 25307
rect 0 24751 577836 25297
rect 0 24741 22777 24751
rect 0 24209 37221 24219
rect 0 23663 577836 24209
rect 0 23653 28389 23663
rect 0 23121 55897 23131
rect 0 22575 577836 23121
rect 0 22565 78897 22575
rect 0 22033 39889 22043
rect 0 21487 577836 22033
rect 0 21477 36301 21487
rect 0 20945 9529 20955
rect 0 20399 577836 20945
rect 0 20389 32345 20399
rect 0 19857 25629 19867
rect 0 19311 577836 19857
rect 0 19301 140629 19311
rect 0 18769 40257 18779
rect 0 18223 577836 18769
rect 0 18213 5941 18223
rect 0 17681 13025 17691
rect 0 17135 577836 17681
rect 0 17125 20201 17135
rect 0 16593 76137 16603
rect 0 16047 577836 16593
rect 0 16037 67673 16047
rect 0 15505 48261 15515
rect 0 14959 577836 15505
rect 0 14949 24617 14959
rect 0 14417 6677 14427
rect 0 13871 577836 14417
rect 0 13861 34185 13871
rect 0 13329 23513 13339
rect 0 12783 577836 13329
rect 0 12773 14405 12783
rect 0 12241 22317 12251
rect 0 11695 577836 12241
rect 0 11685 23605 11695
rect 0 11153 10449 11163
rect 0 10607 577836 11153
rect 0 10597 11553 10607
rect 0 10065 33541 10075
rect 0 9519 577836 10065
rect 0 9509 17165 9519
rect 0 8977 20201 8987
rect 0 8431 577836 8977
rect 0 8421 136949 8431
rect 0 7889 129037 7899
rect 0 7343 577836 7889
rect 0 7333 137685 7343
rect 0 6801 143573 6811
rect 0 6255 577836 6801
rect 0 6245 158937 6255
rect 0 5713 161789 5723
rect 0 5167 577836 5713
rect 0 5157 149369 5167
rect 0 4625 167769 4635
rect 0 4079 577836 4625
rect 0 4069 241645 4079
rect 0 3537 235297 3547
rect 0 2981 577836 3537
rect 0 2138 577836 2459
<< obsli1 >>
rect 38 2159 577953 617457
<< obsm1 >>
rect 38 1980 577965 617488
<< metal2 >>
rect 2356 0 2412 800
rect 9256 0 9312 800
rect 16248 0 16304 800
rect 23240 0 23296 800
rect 30232 0 30288 800
rect 37224 0 37280 800
rect 44216 0 44272 800
rect 51208 0 51264 800
rect 58200 0 58256 800
rect 65192 0 65248 800
rect 72184 0 72240 800
rect 79176 0 79232 800
rect 86168 0 86224 800
rect 93160 0 93216 800
rect 100152 0 100208 800
rect 107144 0 107200 800
rect 114136 0 114192 800
rect 121128 0 121184 800
rect 128120 0 128176 800
rect 135112 0 135168 800
rect 142104 0 142160 800
rect 149004 0 149060 800
rect 155996 0 156052 800
rect 162988 0 163044 800
rect 169980 0 170036 800
rect 176972 0 177028 800
rect 183964 0 184020 800
rect 190956 0 191012 800
rect 197948 0 198004 800
rect 204940 0 204996 800
rect 211932 0 211988 800
rect 218924 0 218980 800
rect 225916 0 225972 800
rect 232908 0 232964 800
rect 239900 0 239956 800
rect 246892 0 246948 800
rect 253884 0 253940 800
rect 260876 0 260932 800
rect 267868 0 267924 800
rect 274860 0 274916 800
rect 281852 0 281908 800
rect 288844 0 288900 800
rect 295744 0 295800 800
rect 302736 0 302792 800
rect 309728 0 309784 800
rect 316720 0 316776 800
rect 323712 0 323768 800
rect 330704 0 330760 800
rect 337696 0 337752 800
rect 344688 0 344744 800
rect 351680 0 351736 800
rect 358672 0 358728 800
rect 365664 0 365720 800
rect 372656 0 372712 800
rect 379648 0 379704 800
rect 386640 0 386696 800
rect 393632 0 393688 800
rect 400624 0 400680 800
rect 407616 0 407672 800
rect 414608 0 414664 800
rect 421600 0 421656 800
rect 428592 0 428648 800
rect 435584 0 435640 800
rect 442484 0 442540 800
rect 449476 0 449532 800
rect 456468 0 456524 800
rect 463460 0 463516 800
rect 470452 0 470508 800
rect 477444 0 477500 800
rect 484436 0 484492 800
rect 491428 0 491484 800
rect 498420 0 498476 800
rect 505412 0 505468 800
rect 512404 0 512460 800
rect 519396 0 519452 800
rect 526388 0 526444 800
rect 533380 0 533436 800
rect 540372 0 540428 800
rect 547364 0 547420 800
rect 554356 0 554412 800
rect 561348 0 561404 800
rect 568340 0 568396 800
rect 575332 0 575388 800
<< obsm2 >>
rect 334 856 577594 617488
rect 334 800 2300 856
rect 2468 800 9200 856
rect 9368 800 16192 856
rect 16360 800 23184 856
rect 23352 800 30176 856
rect 30344 800 37168 856
rect 37336 800 44160 856
rect 44328 800 51152 856
rect 51320 800 58144 856
rect 58312 800 65136 856
rect 65304 800 72128 856
rect 72296 800 79120 856
rect 79288 800 86112 856
rect 86280 800 93104 856
rect 93272 800 100096 856
rect 100264 800 107088 856
rect 107256 800 114080 856
rect 114248 800 121072 856
rect 121240 800 128064 856
rect 128232 800 135056 856
rect 135224 800 142048 856
rect 142216 800 148948 856
rect 149116 800 155940 856
rect 156108 800 162932 856
rect 163100 800 169924 856
rect 170092 800 176916 856
rect 177084 800 183908 856
rect 184076 800 190900 856
rect 191068 800 197892 856
rect 198060 800 204884 856
rect 205052 800 211876 856
rect 212044 800 218868 856
rect 219036 800 225860 856
rect 226028 800 232852 856
rect 233020 800 239844 856
rect 240012 800 246836 856
rect 247004 800 253828 856
rect 253996 800 260820 856
rect 260988 800 267812 856
rect 267980 800 274804 856
rect 274972 800 281796 856
rect 281964 800 288788 856
rect 288956 800 295688 856
rect 295856 800 302680 856
rect 302848 800 309672 856
rect 309840 800 316664 856
rect 316832 800 323656 856
rect 323824 800 330648 856
rect 330816 800 337640 856
rect 337808 800 344632 856
rect 344800 800 351624 856
rect 351792 800 358616 856
rect 358784 800 365608 856
rect 365776 800 372600 856
rect 372768 800 379592 856
rect 379760 800 386584 856
rect 386752 800 393576 856
rect 393744 800 400568 856
rect 400736 800 407560 856
rect 407728 800 414552 856
rect 414720 800 421544 856
rect 421712 800 428536 856
rect 428704 800 435528 856
rect 435696 800 442428 856
rect 442596 800 449420 856
rect 449588 800 456412 856
rect 456580 800 463404 856
rect 463572 800 470396 856
rect 470564 800 477388 856
rect 477556 800 484380 856
rect 484548 800 491372 856
rect 491540 800 498364 856
rect 498532 800 505356 856
rect 505524 800 512348 856
rect 512516 800 519340 856
rect 519508 800 526332 856
rect 526500 800 533324 856
rect 533492 800 540316 856
rect 540484 800 547308 856
rect 547476 800 554300 856
rect 554468 800 561292 856
rect 561460 800 568284 856
rect 568452 800 575276 856
rect 575444 800 577594 856
<< obsm3 >>
rect 971 2143 577417 617473
<< metal4 >>
rect 3142 2128 3462 617488
rect 18502 2128 18822 617488
rect 33862 2128 34182 617488
rect 49222 2128 49542 617488
rect 64582 2128 64902 617488
rect 79942 2128 80262 617488
rect 95302 2128 95622 617488
rect 110662 2128 110982 617488
rect 126022 2128 126342 617488
rect 141382 2128 141702 617488
rect 156742 2128 157062 617488
rect 172102 2128 172422 617488
rect 187462 2128 187782 617488
rect 202822 2128 203142 617488
rect 218182 2128 218502 617488
rect 233542 2128 233862 617488
rect 248902 2128 249222 617488
rect 264262 2128 264582 617488
rect 279622 2128 279942 617488
rect 294982 2128 295302 617488
rect 310342 2128 310662 617488
rect 325702 2128 326022 617488
rect 341062 2128 341382 617488
rect 356422 2128 356742 617488
rect 371782 2128 372102 617488
rect 387142 2128 387462 617488
rect 402502 2128 402822 617488
rect 417862 2128 418182 617488
rect 433222 2128 433542 617488
rect 448582 2128 448902 617488
rect 463942 2128 464262 617488
rect 479302 2128 479622 617488
rect 494662 2128 494982 617488
rect 510022 2128 510342 617488
rect 525382 2128 525702 617488
rect 540742 2128 541062 617488
rect 556102 2128 556422 617488
rect 571462 2128 571782 617488
<< obsm4 >>
rect 3593 2619 18422 611285
rect 18902 2619 33782 611285
rect 34262 2619 49142 611285
rect 49622 2619 64502 611285
rect 64982 2619 79862 611285
rect 80342 2619 95222 611285
rect 95702 2619 110582 611285
rect 111062 2619 125942 611285
rect 126422 2619 141302 611285
rect 141782 2619 156662 611285
rect 157142 2619 172022 611285
rect 172502 2619 187382 611285
rect 187862 2619 202742 611285
rect 203222 2619 218102 611285
rect 218582 2619 233462 611285
rect 233942 2619 248822 611285
rect 249302 2619 264182 611285
rect 264662 2619 279542 611285
rect 280022 2619 294902 611285
rect 295382 2619 310262 611285
rect 310742 2619 325622 611285
rect 326102 2619 340982 611285
rect 341462 2619 356342 611285
rect 356822 2619 371702 611285
rect 372182 2619 387062 611285
rect 387542 2619 402422 611285
rect 402902 2619 417782 611285
rect 418262 2619 433142 611285
rect 433622 2619 448502 611285
rect 448982 2619 463862 611285
rect 464342 2619 479222 611285
rect 479702 2619 494582 611285
rect 495062 2619 509942 611285
rect 510422 2619 525302 611285
rect 525782 2619 540662 611285
rect 541142 2619 556022 611285
rect 556502 2619 561363 611285
<< labels >>
rlabel metal2 s 449476 0 449532 800 6 A[0]
port 1 nsew signal input
rlabel metal2 s 519396 0 519452 800 6 A[10]
port 2 nsew signal input
rlabel metal2 s 526388 0 526444 800 6 A[11]
port 3 nsew signal input
rlabel metal2 s 533380 0 533436 800 6 A[12]
port 4 nsew signal input
rlabel metal2 s 456468 0 456524 800 6 A[1]
port 5 nsew signal input
rlabel metal2 s 463460 0 463516 800 6 A[2]
port 6 nsew signal input
rlabel metal2 s 470452 0 470508 800 6 A[3]
port 7 nsew signal input
rlabel metal2 s 477444 0 477500 800 6 A[4]
port 8 nsew signal input
rlabel metal2 s 484436 0 484492 800 6 A[5]
port 9 nsew signal input
rlabel metal2 s 491428 0 491484 800 6 A[6]
port 10 nsew signal input
rlabel metal2 s 498420 0 498476 800 6 A[7]
port 11 nsew signal input
rlabel metal2 s 505412 0 505468 800 6 A[8]
port 12 nsew signal input
rlabel metal2 s 512404 0 512460 800 6 A[9]
port 13 nsew signal input
rlabel metal2 s 540372 0 540428 800 6 CLK
port 14 nsew signal input
rlabel metal2 s 225916 0 225972 800 6 Di[0]
port 15 nsew signal input
rlabel metal2 s 295744 0 295800 800 6 Di[10]
port 16 nsew signal input
rlabel metal2 s 302736 0 302792 800 6 Di[11]
port 17 nsew signal input
rlabel metal2 s 309728 0 309784 800 6 Di[12]
port 18 nsew signal input
rlabel metal2 s 316720 0 316776 800 6 Di[13]
port 19 nsew signal input
rlabel metal2 s 323712 0 323768 800 6 Di[14]
port 20 nsew signal input
rlabel metal2 s 330704 0 330760 800 6 Di[15]
port 21 nsew signal input
rlabel metal2 s 337696 0 337752 800 6 Di[16]
port 22 nsew signal input
rlabel metal2 s 344688 0 344744 800 6 Di[17]
port 23 nsew signal input
rlabel metal2 s 351680 0 351736 800 6 Di[18]
port 24 nsew signal input
rlabel metal2 s 358672 0 358728 800 6 Di[19]
port 25 nsew signal input
rlabel metal2 s 232908 0 232964 800 6 Di[1]
port 26 nsew signal input
rlabel metal2 s 365664 0 365720 800 6 Di[20]
port 27 nsew signal input
rlabel metal2 s 372656 0 372712 800 6 Di[21]
port 28 nsew signal input
rlabel metal2 s 379648 0 379704 800 6 Di[22]
port 29 nsew signal input
rlabel metal2 s 386640 0 386696 800 6 Di[23]
port 30 nsew signal input
rlabel metal2 s 393632 0 393688 800 6 Di[24]
port 31 nsew signal input
rlabel metal2 s 400624 0 400680 800 6 Di[25]
port 32 nsew signal input
rlabel metal2 s 407616 0 407672 800 6 Di[26]
port 33 nsew signal input
rlabel metal2 s 414608 0 414664 800 6 Di[27]
port 34 nsew signal input
rlabel metal2 s 421600 0 421656 800 6 Di[28]
port 35 nsew signal input
rlabel metal2 s 428592 0 428648 800 6 Di[29]
port 36 nsew signal input
rlabel metal2 s 239900 0 239956 800 6 Di[2]
port 37 nsew signal input
rlabel metal2 s 435584 0 435640 800 6 Di[30]
port 38 nsew signal input
rlabel metal2 s 442484 0 442540 800 6 Di[31]
port 39 nsew signal input
rlabel metal2 s 246892 0 246948 800 6 Di[3]
port 40 nsew signal input
rlabel metal2 s 253884 0 253940 800 6 Di[4]
port 41 nsew signal input
rlabel metal2 s 260876 0 260932 800 6 Di[5]
port 42 nsew signal input
rlabel metal2 s 267868 0 267924 800 6 Di[6]
port 43 nsew signal input
rlabel metal2 s 274860 0 274916 800 6 Di[7]
port 44 nsew signal input
rlabel metal2 s 281852 0 281908 800 6 Di[8]
port 45 nsew signal input
rlabel metal2 s 288844 0 288900 800 6 Di[9]
port 46 nsew signal input
rlabel metal2 s 2356 0 2412 800 6 Do[0]
port 47 nsew signal output
rlabel metal2 s 72184 0 72240 800 6 Do[10]
port 48 nsew signal output
rlabel metal2 s 79176 0 79232 800 6 Do[11]
port 49 nsew signal output
rlabel metal2 s 86168 0 86224 800 6 Do[12]
port 50 nsew signal output
rlabel metal2 s 93160 0 93216 800 6 Do[13]
port 51 nsew signal output
rlabel metal2 s 100152 0 100208 800 6 Do[14]
port 52 nsew signal output
rlabel metal2 s 107144 0 107200 800 6 Do[15]
port 53 nsew signal output
rlabel metal2 s 114136 0 114192 800 6 Do[16]
port 54 nsew signal output
rlabel metal2 s 121128 0 121184 800 6 Do[17]
port 55 nsew signal output
rlabel metal2 s 128120 0 128176 800 6 Do[18]
port 56 nsew signal output
rlabel metal2 s 135112 0 135168 800 6 Do[19]
port 57 nsew signal output
rlabel metal2 s 9256 0 9312 800 6 Do[1]
port 58 nsew signal output
rlabel metal2 s 142104 0 142160 800 6 Do[20]
port 59 nsew signal output
rlabel metal2 s 149004 0 149060 800 6 Do[21]
port 60 nsew signal output
rlabel metal2 s 155996 0 156052 800 6 Do[22]
port 61 nsew signal output
rlabel metal2 s 162988 0 163044 800 6 Do[23]
port 62 nsew signal output
rlabel metal2 s 169980 0 170036 800 6 Do[24]
port 63 nsew signal output
rlabel metal2 s 176972 0 177028 800 6 Do[25]
port 64 nsew signal output
rlabel metal2 s 183964 0 184020 800 6 Do[26]
port 65 nsew signal output
rlabel metal2 s 190956 0 191012 800 6 Do[27]
port 66 nsew signal output
rlabel metal2 s 197948 0 198004 800 6 Do[28]
port 67 nsew signal output
rlabel metal2 s 204940 0 204996 800 6 Do[29]
port 68 nsew signal output
rlabel metal2 s 16248 0 16304 800 6 Do[2]
port 69 nsew signal output
rlabel metal2 s 211932 0 211988 800 6 Do[30]
port 70 nsew signal output
rlabel metal2 s 218924 0 218980 800 6 Do[31]
port 71 nsew signal output
rlabel metal2 s 23240 0 23296 800 6 Do[3]
port 72 nsew signal output
rlabel metal2 s 30232 0 30288 800 6 Do[4]
port 73 nsew signal output
rlabel metal2 s 37224 0 37280 800 6 Do[5]
port 74 nsew signal output
rlabel metal2 s 44216 0 44272 800 6 Do[6]
port 75 nsew signal output
rlabel metal2 s 51208 0 51264 800 6 Do[7]
port 76 nsew signal output
rlabel metal2 s 58200 0 58256 800 6 Do[8]
port 77 nsew signal output
rlabel metal2 s 65192 0 65248 800 6 Do[9]
port 78 nsew signal output
rlabel metal2 s 575332 0 575388 800 6 EN
port 79 nsew signal input
rlabel metal2 s 547364 0 547420 800 6 WE[0]
port 80 nsew signal input
rlabel metal2 s 554356 0 554412 800 6 WE[1]
port 81 nsew signal input
rlabel metal2 s 561348 0 561404 800 6 WE[2]
port 82 nsew signal input
rlabel metal2 s 568340 0 568396 800 6 WE[3]
port 83 nsew signal input
rlabel metal4 s 556102 2128 556422 617488 6 VPWR
port 84 nsew power bidirectional
rlabel metal4 s 525382 2128 525702 617488 6 VPWR
port 85 nsew power bidirectional
rlabel metal4 s 494662 2128 494982 617488 6 VPWR
port 86 nsew power bidirectional
rlabel metal4 s 463942 2128 464262 617488 6 VPWR
port 87 nsew power bidirectional
rlabel metal4 s 433222 2128 433542 617488 6 VPWR
port 88 nsew power bidirectional
rlabel metal4 s 402502 2128 402822 617488 6 VPWR
port 89 nsew power bidirectional
rlabel metal4 s 371782 2128 372102 617488 6 VPWR
port 90 nsew power bidirectional
rlabel metal4 s 341062 2128 341382 617488 6 VPWR
port 91 nsew power bidirectional
rlabel metal4 s 310342 2128 310662 617488 6 VPWR
port 92 nsew power bidirectional
rlabel metal4 s 279622 2128 279942 617488 6 VPWR
port 93 nsew power bidirectional
rlabel metal4 s 248902 2128 249222 617488 6 VPWR
port 94 nsew power bidirectional
rlabel metal4 s 218182 2128 218502 617488 6 VPWR
port 95 nsew power bidirectional
rlabel metal4 s 187462 2128 187782 617488 6 VPWR
port 96 nsew power bidirectional
rlabel metal4 s 156742 2128 157062 617488 6 VPWR
port 97 nsew power bidirectional
rlabel metal4 s 126022 2128 126342 617488 6 VPWR
port 98 nsew power bidirectional
rlabel metal4 s 95302 2128 95622 617488 6 VPWR
port 99 nsew power bidirectional
rlabel metal4 s 64582 2128 64902 617488 6 VPWR
port 100 nsew power bidirectional
rlabel metal4 s 33862 2128 34182 617488 6 VPWR
port 101 nsew power bidirectional
rlabel metal4 s 3142 2128 3462 617488 6 VPWR
port 102 nsew power bidirectional
rlabel metal4 s 571462 2128 571782 617488 6 VGND
port 103 nsew ground bidirectional
rlabel metal4 s 540742 2128 541062 617488 6 VGND
port 104 nsew ground bidirectional
rlabel metal4 s 510022 2128 510342 617488 6 VGND
port 105 nsew ground bidirectional
rlabel metal4 s 479302 2128 479622 617488 6 VGND
port 106 nsew ground bidirectional
rlabel metal4 s 448582 2128 448902 617488 6 VGND
port 107 nsew ground bidirectional
rlabel metal4 s 417862 2128 418182 617488 6 VGND
port 108 nsew ground bidirectional
rlabel metal4 s 387142 2128 387462 617488 6 VGND
port 109 nsew ground bidirectional
rlabel metal4 s 356422 2128 356742 617488 6 VGND
port 110 nsew ground bidirectional
rlabel metal4 s 325702 2128 326022 617488 6 VGND
port 111 nsew ground bidirectional
rlabel metal4 s 294982 2128 295302 617488 6 VGND
port 112 nsew ground bidirectional
rlabel metal4 s 264262 2128 264582 617488 6 VGND
port 113 nsew ground bidirectional
rlabel metal4 s 233542 2128 233862 617488 6 VGND
port 114 nsew ground bidirectional
rlabel metal4 s 202822 2128 203142 617488 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 172102 2128 172422 617488 6 VGND
port 116 nsew ground bidirectional
rlabel metal4 s 141382 2128 141702 617488 6 VGND
port 117 nsew ground bidirectional
rlabel metal4 s 110662 2128 110982 617488 6 VGND
port 118 nsew ground bidirectional
rlabel metal4 s 79942 2128 80262 617488 6 VGND
port 119 nsew ground bidirectional
rlabel metal4 s 49222 2128 49542 617488 6 VGND
port 120 nsew ground bidirectional
rlabel metal4 s 18502 2128 18822 617488 6 VGND
port 121 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 577965 617488
string LEFview TRUE
string GDS_FILE /project/openlane/RAM_6Kx32/runs/RAM_6Kx32/results/magic/RAM_6Kx32.gds
string GDS_END 1337535352
string GDS_START 226610
<< end >>

