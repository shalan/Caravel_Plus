VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM_6Kx32
  CLASS BLOCK ;
  FOREIGN RAM_6Kx32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2889.825 BY 3087.870 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.380 0.000 2247.660 4.000 ;
    END
  END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2596.980 0.000 2597.260 4.000 ;
    END
  END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2631.940 0.000 2632.220 4.000 ;
    END
  END A[11]
  PIN A[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2666.900 0.000 2667.180 4.000 ;
    END
  END A[12]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.340 0.000 2282.620 4.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2317.300 0.000 2317.580 4.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2352.260 0.000 2352.540 4.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2387.220 0.000 2387.500 4.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.180 0.000 2422.460 4.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2457.140 0.000 2457.420 4.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2492.100 0.000 2492.380 4.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.060 0.000 2527.340 4.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.020 0.000 2562.300 4.000 ;
    END
  END A[9]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2701.860 0.000 2702.140 4.000 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.580 0.000 1129.860 4.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.720 0.000 1479.000 4.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.680 0.000 1513.960 4.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.640 0.000 1548.920 4.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.600 0.000 1583.880 4.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.560 0.000 1618.840 4.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.520 0.000 1653.800 4.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.480 0.000 1688.760 4.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.440 0.000 1723.720 4.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.400 0.000 1758.680 4.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.360 0.000 1793.640 4.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.540 0.000 1164.820 4.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.320 0.000 1828.600 4.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.280 0.000 1863.560 4.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.240 0.000 1898.520 4.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.200 0.000 1933.480 4.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1968.160 0.000 1968.440 4.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.120 0.000 2003.400 4.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.080 0.000 2038.360 4.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.040 0.000 2073.320 4.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.000 0.000 2108.280 4.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.960 0.000 2143.240 4.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.500 0.000 1199.780 4.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.920 0.000 2178.200 4.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.420 0.000 2212.700 4.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.460 0.000 1234.740 4.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.420 0.000 1269.700 4.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.380 0.000 1304.660 4.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.340 0.000 1339.620 4.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.300 0.000 1374.580 4.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.260 0.000 1409.540 4.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.220 0.000 1444.500 4.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.780 0.000 12.060 4.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.920 0.000 361.200 4.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.880 0.000 396.160 4.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.840 0.000 431.120 4.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.800 0.000 466.080 4.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.760 0.000 501.040 4.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.720 0.000 536.000 4.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.680 0.000 570.960 4.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.640 0.000 605.920 4.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.600 0.000 640.880 4.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.560 0.000 675.840 4.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.280 0.000 46.560 4.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.520 0.000 710.800 4.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.020 0.000 745.300 4.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.980 0.000 780.260 4.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.940 0.000 815.220 4.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.900 0.000 850.180 4.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.860 0.000 885.140 4.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.820 0.000 920.100 4.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.780 0.000 955.060 4.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.740 0.000 990.020 4.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.700 0.000 1024.980 4.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.240 0.000 81.520 4.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.660 0.000 1059.940 4.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.620 0.000 1094.900 4.000 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.200 0.000 116.480 4.000 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.160 0.000 151.440 4.000 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.120 0.000 186.400 4.000 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.080 0.000 221.360 4.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.040 0.000 256.320 4.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.000 0.000 291.280 4.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.960 0.000 326.240 4.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2876.660 0.000 2876.940 4.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2736.820 0.000 2737.100 4.000 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2771.780 0.000 2772.060 4.000 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2806.740 0.000 2807.020 4.000 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2841.700 0.000 2841.980 4.000 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2780.510 10.640 2782.110 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2626.910 10.640 2628.510 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2473.310 10.640 2474.910 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2319.710 10.640 2321.310 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2166.110 10.640 2167.710 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2012.510 10.640 2014.110 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1858.910 10.640 1860.510 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1705.310 10.640 1706.910 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1551.710 10.640 1553.310 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1398.110 10.640 1399.710 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1244.510 10.640 1246.110 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1090.910 10.640 1092.510 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 937.310 10.640 938.910 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 783.710 10.640 785.310 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 630.110 10.640 631.710 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 476.510 10.640 478.110 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 322.910 10.640 324.510 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 169.310 10.640 170.910 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.710 10.640 17.310 3087.440 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2857.310 10.640 2858.910 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2703.710 10.640 2705.310 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2550.110 10.640 2551.710 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2396.510 10.640 2398.110 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2242.910 10.640 2244.510 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2089.310 10.640 2090.910 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1935.710 10.640 1937.310 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1782.110 10.640 1783.710 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1628.510 10.640 1630.110 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1474.910 10.640 1476.510 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1321.310 10.640 1322.910 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1167.710 10.640 1169.310 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1014.110 10.640 1015.710 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 860.510 10.640 862.110 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 706.910 10.640 708.510 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 553.310 10.640 554.910 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 399.710 10.640 401.310 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.110 10.640 247.710 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 92.510 10.640 94.110 3087.440 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.000 3083.065 1.760 3085.895 ;
        RECT 0.000 3077.625 1.760 3080.455 ;
        RECT 0.000 3072.185 1.760 3075.015 ;
        RECT 0.000 3066.745 1.760 3069.575 ;
        RECT 0.000 3061.305 1.760 3064.135 ;
        RECT 0.000 3055.865 1.760 3058.695 ;
        RECT 0.000 3050.425 1.760 3053.255 ;
        RECT 0.000 3044.985 1.760 3047.815 ;
        RECT 0.000 3039.545 1.760 3042.375 ;
        RECT 0.000 3034.105 1.760 3036.935 ;
        RECT 0.000 3028.665 1.760 3031.495 ;
        RECT 0.000 3023.225 1.760 3026.055 ;
        RECT 0.000 3019.390 1.760 3020.615 ;
        RECT 0.000 3019.010 33.040 3019.390 ;
        RECT 0.000 3017.785 25.680 3019.010 ;
        RECT 0.000 3013.950 1.760 3015.175 ;
        RECT 0.000 3013.570 394.600 3013.950 ;
        RECT 0.000 3012.345 51.900 3013.570 ;
        RECT 0.000 3006.905 1.760 3009.735 ;
        RECT 0.000 3001.465 1.760 3004.295 ;
        RECT 0.000 2996.025 1.760 2998.855 ;
        RECT 0.000 2990.585 1.760 2993.415 ;
        RECT 0.000 2986.750 1.760 2987.975 ;
        RECT 0.000 2985.145 14.180 2986.750 ;
        RECT 0.000 2979.705 1.760 2982.535 ;
        RECT 0.000 2974.265 1.760 2977.095 ;
        RECT 0.000 2968.825 1.760 2971.655 ;
        RECT 0.000 2963.385 1.760 2966.215 ;
        RECT 0.000 2957.945 1.760 2960.775 ;
        RECT 0.000 2952.505 1.760 2955.335 ;
        RECT 0.000 2947.065 1.760 2949.895 ;
        RECT 0.000 2941.625 1.760 2944.455 ;
        RECT 0.000 2936.185 1.760 2939.015 ;
        RECT 0.000 2930.745 1.760 2933.575 ;
        RECT 0.000 2928.085 2.565 2928.135 ;
        RECT 0.000 2926.910 9.120 2928.085 ;
        RECT 0.000 2926.530 33.040 2926.910 ;
        RECT 0.000 2925.305 1.760 2926.530 ;
        RECT 0.000 2919.865 1.760 2922.695 ;
        RECT 0.000 2914.425 1.760 2917.255 ;
        RECT 0.000 2908.985 1.760 2911.815 ;
        RECT 0.000 2905.150 9.120 2906.375 ;
        RECT 0.000 2904.770 252.000 2905.150 ;
        RECT 0.000 2903.545 1.760 2904.770 ;
        RECT 0.000 2898.105 1.760 2900.935 ;
        RECT 0.000 2894.270 9.120 2895.495 ;
        RECT 0.000 2893.890 231.300 2894.270 ;
        RECT 0.000 2892.715 19.700 2893.890 ;
        RECT 0.000 2892.665 2.565 2892.715 ;
        RECT 0.000 2888.830 9.120 2890.055 ;
        RECT 0.000 2888.450 238.200 2888.830 ;
        RECT 0.000 2887.225 1.760 2888.450 ;
        RECT 0.000 2881.785 1.760 2884.615 ;
        RECT 0.000 2876.345 1.760 2879.175 ;
        RECT 0.000 2870.905 1.760 2873.735 ;
        RECT 0.000 2865.465 1.760 2868.295 ;
        RECT 0.000 2860.025 1.760 2862.855 ;
        RECT 0.000 2854.585 1.760 2857.415 ;
        RECT 0.000 2849.145 1.760 2851.975 ;
        RECT 0.000 2843.705 1.760 2846.535 ;
        RECT 0.000 2838.265 1.760 2841.095 ;
        RECT 0.000 2834.430 10.040 2835.655 ;
        RECT 0.000 2834.050 213.360 2834.430 ;
        RECT 0.000 2832.825 20.620 2834.050 ;
        RECT 0.000 2827.385 1.760 2830.215 ;
        RECT 0.000 2821.945 1.760 2824.775 ;
        RECT 0.000 2816.505 1.760 2819.335 ;
        RECT 0.000 2811.065 1.760 2813.895 ;
        RECT 0.000 2805.625 1.760 2808.455 ;
        RECT 0.000 2800.185 1.760 2803.015 ;
        RECT 0.000 2794.745 1.760 2797.575 ;
        RECT 0.000 2790.910 1.760 2792.135 ;
        RECT 0.000 2790.530 10.500 2790.910 ;
        RECT 0.000 2789.355 10.040 2790.530 ;
        RECT 0.000 2789.305 2.565 2789.355 ;
        RECT 0.000 2783.865 1.760 2786.695 ;
        RECT 0.000 2778.425 1.760 2781.255 ;
        RECT 0.000 2772.985 1.760 2775.815 ;
        RECT 0.000 2767.545 1.760 2770.375 ;
        RECT 0.000 2762.105 1.760 2764.935 ;
        RECT 0.000 2756.665 1.760 2759.495 ;
        RECT 0.000 2751.225 1.760 2754.055 ;
        RECT 0.000 2745.785 1.760 2748.615 ;
        RECT 0.000 2741.950 14.180 2743.175 ;
        RECT 0.000 2741.570 272.700 2741.950 ;
        RECT 0.000 2740.345 27.060 2741.570 ;
        RECT 0.000 2736.510 5.900 2737.735 ;
        RECT 0.000 2736.130 31.200 2736.510 ;
        RECT 0.000 2734.955 27.980 2736.130 ;
        RECT 0.000 2734.905 2.565 2734.955 ;
        RECT 0.000 2729.465 1.760 2732.295 ;
        RECT 0.000 2725.630 1.760 2726.855 ;
        RECT 0.000 2725.250 112.160 2725.630 ;
        RECT 0.000 2724.025 16.020 2725.250 ;
        RECT 0.000 2720.190 10.040 2721.415 ;
        RECT 0.000 2719.810 15.560 2720.190 ;
        RECT 0.000 2718.585 1.760 2719.810 ;
        RECT 0.000 2713.145 1.760 2715.975 ;
        RECT 0.000 2707.705 1.760 2710.535 ;
        RECT 0.000 2702.265 1.760 2705.095 ;
        RECT 0.000 2696.825 1.760 2699.655 ;
        RECT 0.000 2691.385 1.760 2694.215 ;
        RECT 0.000 2685.945 1.760 2688.775 ;
        RECT 0.000 2680.505 1.760 2683.335 ;
        RECT 0.000 2675.065 1.760 2677.895 ;
        RECT 0.000 2669.625 1.760 2672.455 ;
        RECT 0.000 2664.185 1.760 2667.015 ;
        RECT 0.000 2658.745 1.760 2661.575 ;
        RECT 0.000 2653.305 1.760 2656.135 ;
        RECT 0.000 2647.865 1.760 2650.695 ;
        RECT 0.000 2644.030 9.120 2645.255 ;
        RECT 0.000 2643.650 13.720 2644.030 ;
        RECT 0.000 2642.425 1.760 2643.650 ;
        RECT 0.000 2636.985 1.760 2639.815 ;
        RECT 0.000 2634.325 2.565 2634.375 ;
        RECT 0.000 2633.150 42.240 2634.325 ;
        RECT 0.000 2632.770 104.340 2633.150 ;
        RECT 0.000 2631.545 1.760 2632.770 ;
        RECT 0.000 2627.710 9.120 2628.935 ;
        RECT 0.000 2627.330 70.300 2627.710 ;
        RECT 0.000 2626.105 15.100 2627.330 ;
        RECT 0.000 2620.665 1.760 2623.495 ;
        RECT 0.000 2616.830 10.040 2618.055 ;
        RECT 0.000 2616.450 125.500 2616.830 ;
        RECT 0.000 2615.225 1.760 2616.450 ;
        RECT 0.000 2611.010 14.180 2612.615 ;
        RECT 0.000 2609.785 1.760 2611.010 ;
        RECT 0.000 2605.950 9.120 2607.175 ;
        RECT 0.000 2605.570 124.120 2605.950 ;
        RECT 0.000 2604.345 1.760 2605.570 ;
        RECT 0.000 2598.905 1.760 2601.735 ;
        RECT 0.000 2593.465 1.760 2596.295 ;
        RECT 0.000 2588.025 1.760 2590.855 ;
        RECT 0.000 2584.190 1.760 2585.415 ;
        RECT 0.000 2582.635 9.120 2584.190 ;
        RECT 0.000 2582.585 2.565 2582.635 ;
        RECT 0.000 2578.750 1.760 2579.975 ;
        RECT 0.000 2578.370 448.420 2578.750 ;
        RECT 0.000 2577.145 26.600 2578.370 ;
        RECT 0.000 2571.705 1.760 2574.535 ;
        RECT 0.000 2566.265 1.760 2569.095 ;
        RECT 0.000 2560.825 1.760 2563.655 ;
        RECT 0.000 2555.385 1.760 2558.215 ;
        RECT 0.000 2551.550 1.760 2552.775 ;
        RECT 0.000 2551.170 97.440 2551.550 ;
        RECT 0.000 2549.995 27.980 2551.170 ;
        RECT 0.000 2549.945 9.925 2549.995 ;
        RECT 0.000 2544.505 1.760 2547.335 ;
        RECT 0.000 2540.670 1.760 2541.895 ;
        RECT 0.000 2540.290 67.080 2540.670 ;
        RECT 0.000 2539.065 9.120 2540.290 ;
        RECT 0.000 2533.625 1.760 2536.455 ;
        RECT 0.000 2528.185 1.760 2531.015 ;
        RECT 0.000 2522.745 14.180 2525.575 ;
        RECT 0.000 2517.305 1.760 2520.135 ;
        RECT 0.000 2513.470 10.040 2514.695 ;
        RECT 0.000 2513.090 235.440 2513.470 ;
        RECT 0.000 2511.915 10.500 2513.090 ;
        RECT 0.000 2511.865 2.565 2511.915 ;
        RECT 0.000 2508.030 15.100 2509.255 ;
        RECT 0.000 2507.650 168.280 2508.030 ;
        RECT 0.000 2506.425 14.180 2507.650 ;
        RECT 0.000 2500.985 1.760 2503.815 ;
        RECT 0.000 2497.150 1.760 2498.375 ;
        RECT 0.000 2496.770 29.820 2497.150 ;
        RECT 0.000 2495.545 16.480 2496.770 ;
        RECT 0.000 2491.710 14.180 2492.935 ;
        RECT 0.000 2491.330 44.080 2491.710 ;
        RECT 0.000 2490.105 1.760 2491.330 ;
        RECT 0.000 2486.270 10.040 2487.495 ;
        RECT 0.000 2485.890 78.120 2486.270 ;
        RECT 0.000 2484.665 1.760 2485.890 ;
        RECT 0.000 2480.830 9.120 2482.055 ;
        RECT 0.000 2480.450 110.320 2480.830 ;
        RECT 0.000 2479.225 1.760 2480.450 ;
        RECT 0.000 2476.565 2.565 2476.615 ;
        RECT 0.000 2475.390 14.180 2476.565 ;
        RECT 0.000 2475.010 19.240 2475.390 ;
        RECT 0.000 2473.785 5.900 2475.010 ;
        RECT 0.000 2469.950 1.760 2471.175 ;
        RECT 0.000 2469.570 566.180 2469.950 ;
        RECT 0.000 2468.395 15.560 2469.570 ;
        RECT 0.000 2468.345 9.925 2468.395 ;
        RECT 0.000 2464.510 9.120 2465.735 ;
        RECT 0.000 2464.130 47.300 2464.510 ;
        RECT 0.000 2462.905 1.760 2464.130 ;
        RECT 0.000 2457.465 1.760 2460.295 ;
        RECT 0.000 2453.630 1.760 2454.855 ;
        RECT 0.000 2453.250 78.580 2453.630 ;
        RECT 0.000 2452.075 9.120 2453.250 ;
        RECT 0.000 2452.025 2.565 2452.075 ;
        RECT 0.000 2446.585 1.760 2449.415 ;
        RECT 0.000 2441.145 1.760 2443.975 ;
        RECT 0.000 2435.705 1.760 2438.535 ;
        RECT 0.000 2430.265 1.760 2433.095 ;
        RECT 0.000 2424.825 1.760 2427.655 ;
        RECT 0.000 2419.385 1.760 2422.215 ;
        RECT 0.000 2416.725 2.565 2416.775 ;
        RECT 0.000 2415.550 9.120 2416.725 ;
        RECT 0.000 2415.170 55.580 2415.550 ;
        RECT 0.000 2413.945 1.760 2415.170 ;
        RECT 0.000 2410.110 19.240 2411.335 ;
        RECT 0.000 2409.730 56.040 2410.110 ;
        RECT 0.000 2408.505 1.760 2409.730 ;
        RECT 0.000 2404.670 10.040 2405.895 ;
        RECT 0.000 2404.290 280.060 2404.670 ;
        RECT 0.000 2403.065 27.980 2404.290 ;
        RECT 0.000 2399.230 14.180 2400.455 ;
        RECT 0.000 2398.850 140.220 2399.230 ;
        RECT 0.000 2397.625 1.760 2398.850 ;
        RECT 0.000 2394.965 2.565 2395.015 ;
        RECT 0.000 2393.790 9.120 2394.965 ;
        RECT 0.000 2393.410 113.080 2393.790 ;
        RECT 0.000 2392.185 1.760 2393.410 ;
        RECT 0.000 2388.350 42.240 2389.575 ;
        RECT 0.000 2387.970 55.120 2388.350 ;
        RECT 0.000 2386.745 1.760 2387.970 ;
        RECT 0.000 2381.305 1.760 2384.135 ;
        RECT 0.000 2375.865 1.760 2378.695 ;
        RECT 0.000 2372.030 1.760 2373.255 ;
        RECT 0.000 2370.425 17.400 2372.030 ;
        RECT 0.000 2366.590 1.760 2367.815 ;
        RECT 0.000 2366.210 42.240 2366.590 ;
        RECT 0.000 2364.985 27.980 2366.210 ;
        RECT 0.000 2362.325 2.565 2362.375 ;
        RECT 0.000 2361.150 27.520 2362.325 ;
        RECT 0.000 2360.770 57.880 2361.150 ;
        RECT 0.000 2359.545 1.760 2360.770 ;
        RECT 0.000 2355.710 1.760 2356.935 ;
        RECT 0.000 2354.105 14.180 2355.710 ;
        RECT 0.000 2350.270 14.180 2351.495 ;
        RECT 0.000 2349.890 75.360 2350.270 ;
        RECT 0.000 2348.665 13.260 2349.890 ;
        RECT 0.000 2343.225 1.760 2346.055 ;
        RECT 0.000 2337.785 1.760 2340.615 ;
        RECT 0.000 2332.345 1.760 2335.175 ;
        RECT 0.000 2326.905 1.760 2329.735 ;
        RECT 0.000 2321.465 1.760 2324.295 ;
        RECT 0.000 2316.025 1.760 2318.855 ;
        RECT 0.000 2310.585 1.760 2313.415 ;
        RECT 0.000 2305.145 1.760 2307.975 ;
        RECT 0.000 2299.705 1.760 2302.535 ;
        RECT 0.000 2295.870 16.020 2297.095 ;
        RECT 0.000 2295.490 277.300 2295.870 ;
        RECT 0.000 2294.265 1.760 2295.490 ;
        RECT 0.000 2291.605 2.565 2291.655 ;
        RECT 0.000 2290.430 22.460 2291.605 ;
        RECT 0.000 2290.050 352.740 2290.430 ;
        RECT 0.000 2288.825 1.760 2290.050 ;
        RECT 0.000 2283.385 1.760 2286.215 ;
        RECT 0.000 2277.945 1.760 2280.775 ;
        RECT 0.000 2274.110 1.760 2275.335 ;
        RECT 0.000 2272.505 18.320 2274.110 ;
        RECT 0.000 2268.670 14.180 2269.895 ;
        RECT 0.000 2268.290 111.700 2268.670 ;
        RECT 0.000 2267.065 1.760 2268.290 ;
        RECT 0.000 2261.625 1.760 2264.455 ;
        RECT 0.000 2257.790 14.180 2259.015 ;
        RECT 0.000 2257.410 84.100 2257.790 ;
        RECT 0.000 2256.185 1.760 2257.410 ;
        RECT 0.000 2252.350 1.760 2253.575 ;
        RECT 0.000 2251.970 210.600 2252.350 ;
        RECT 0.000 2250.795 10.040 2251.970 ;
        RECT 0.000 2250.745 2.565 2250.795 ;
        RECT 0.000 2246.910 1.760 2248.135 ;
        RECT 0.000 2246.530 96.980 2246.910 ;
        RECT 0.000 2245.355 10.500 2246.530 ;
        RECT 0.000 2245.305 2.565 2245.355 ;
        RECT 0.000 2239.865 1.760 2242.695 ;
        RECT 0.000 2234.425 1.760 2237.255 ;
        RECT 0.000 2230.590 9.120 2231.815 ;
        RECT 0.000 2230.210 212.900 2230.590 ;
        RECT 0.000 2228.985 1.760 2230.210 ;
        RECT 0.000 2223.545 1.760 2226.375 ;
        RECT 0.000 2218.105 1.760 2220.935 ;
        RECT 0.000 2212.665 1.760 2215.495 ;
        RECT 0.000 2207.225 1.760 2210.055 ;
        RECT 0.000 2203.390 1.760 2204.615 ;
        RECT 0.000 2203.010 34.420 2203.390 ;
        RECT 0.000 2201.785 9.120 2203.010 ;
        RECT 0.000 2196.345 1.760 2199.175 ;
        RECT 0.000 2190.905 1.760 2193.735 ;
        RECT 0.000 2188.245 2.565 2188.295 ;
        RECT 0.000 2187.070 9.120 2188.245 ;
        RECT 0.000 2186.690 27.980 2187.070 ;
        RECT 0.000 2185.465 1.760 2186.690 ;
        RECT 0.000 2180.025 1.760 2182.855 ;
        RECT 0.000 2174.585 1.760 2177.415 ;
        RECT 0.000 2169.145 1.760 2171.975 ;
        RECT 0.000 2165.310 1.760 2166.535 ;
        RECT 0.000 2164.930 182.080 2165.310 ;
        RECT 0.000 2163.705 17.400 2164.930 ;
        RECT 0.000 2158.265 1.760 2161.095 ;
        RECT 0.000 2155.605 2.565 2155.655 ;
        RECT 0.000 2154.430 9.120 2155.605 ;
        RECT 0.000 2154.050 19.700 2154.430 ;
        RECT 0.000 2152.825 1.760 2154.050 ;
        RECT 0.000 2148.990 1.760 2150.215 ;
        RECT 0.000 2148.610 64.320 2148.990 ;
        RECT 0.000 2147.435 27.980 2148.610 ;
        RECT 0.000 2147.385 14.985 2147.435 ;
        RECT 0.000 2144.725 2.565 2144.775 ;
        RECT 0.000 2143.550 9.120 2144.725 ;
        RECT 0.000 2143.170 332.500 2143.550 ;
        RECT 0.000 2141.945 1.760 2143.170 ;
        RECT 0.000 2136.505 1.760 2139.335 ;
        RECT 0.000 2132.670 1.760 2133.895 ;
        RECT 0.000 2132.290 42.240 2132.670 ;
        RECT 0.000 2131.065 10.040 2132.290 ;
        RECT 0.000 2127.230 1.760 2128.455 ;
        RECT 0.000 2126.850 30.740 2127.230 ;
        RECT 0.000 2125.625 18.320 2126.850 ;
        RECT 0.000 2120.185 1.760 2123.015 ;
        RECT 0.000 2114.745 1.760 2117.575 ;
        RECT 0.000 2109.305 1.760 2112.135 ;
        RECT 0.000 2103.865 1.760 2106.695 ;
        RECT 0.000 2100.030 12.340 2101.255 ;
        RECT 0.000 2099.650 29.360 2100.030 ;
        RECT 0.000 2098.425 1.760 2099.650 ;
        RECT 0.000 2095.765 2.565 2095.815 ;
        RECT 0.000 2094.210 9.120 2095.765 ;
        RECT 0.000 2092.985 1.760 2094.210 ;
        RECT 0.000 2087.545 1.760 2090.375 ;
        RECT 0.000 2083.330 16.020 2084.935 ;
        RECT 0.000 2082.105 10.960 2083.330 ;
        RECT 0.000 2076.665 1.760 2079.495 ;
        RECT 0.000 2072.450 14.180 2074.055 ;
        RECT 0.000 2071.225 1.760 2072.450 ;
        RECT 0.000 2065.785 14.180 2068.615 ;
        RECT 0.000 2060.345 1.760 2063.175 ;
        RECT 0.000 2054.905 1.760 2057.735 ;
        RECT 0.000 2049.465 1.760 2052.295 ;
        RECT 0.000 2044.025 1.760 2046.855 ;
        RECT 0.000 2038.585 1.760 2041.415 ;
        RECT 0.000 2033.145 1.760 2035.975 ;
        RECT 0.000 2027.705 1.760 2030.535 ;
        RECT 0.000 2022.265 1.760 2025.095 ;
        RECT 0.000 2016.825 1.760 2019.655 ;
        RECT 0.000 2011.385 1.760 2014.215 ;
        RECT 0.000 2005.945 1.760 2008.775 ;
        RECT 0.000 2002.110 1.760 2003.335 ;
        RECT 0.000 2001.730 50.520 2002.110 ;
        RECT 0.000 2000.555 19.700 2001.730 ;
        RECT 0.000 2000.505 2.565 2000.555 ;
        RECT 0.000 1995.065 1.760 1997.895 ;
        RECT 0.000 1989.625 1.760 1992.455 ;
        RECT 0.000 1984.185 1.760 1987.015 ;
        RECT 0.000 1978.745 1.760 1981.575 ;
        RECT 0.000 1973.305 1.760 1976.135 ;
        RECT 0.000 1967.865 1.760 1970.695 ;
        RECT 0.000 1962.425 1.760 1965.255 ;
        RECT 0.000 1956.985 1.760 1959.815 ;
        RECT 0.000 1951.545 1.760 1954.375 ;
        RECT 0.000 1946.105 1.760 1948.935 ;
        RECT 0.000 1940.665 1.760 1943.495 ;
        RECT 0.000 1936.830 9.120 1938.055 ;
        RECT 0.000 1936.450 463.140 1936.830 ;
        RECT 0.000 1935.225 1.760 1936.450 ;
        RECT 0.000 1929.785 1.760 1932.615 ;
        RECT 0.000 1927.125 2.565 1927.175 ;
        RECT 0.000 1925.950 9.120 1927.125 ;
        RECT 0.000 1925.570 250.160 1925.950 ;
        RECT 0.000 1924.345 1.760 1925.570 ;
        RECT 0.000 1918.905 1.760 1921.735 ;
        RECT 0.000 1913.465 1.760 1916.295 ;
        RECT 0.000 1908.025 1.760 1910.855 ;
        RECT 0.000 1904.190 1.760 1905.415 ;
        RECT 0.000 1903.810 156.320 1904.190 ;
        RECT 0.000 1902.635 23.840 1903.810 ;
        RECT 0.000 1902.585 2.565 1902.635 ;
        RECT 0.000 1897.145 1.760 1899.975 ;
        RECT 0.000 1893.310 1.760 1894.535 ;
        RECT 0.000 1892.930 81.800 1893.310 ;
        RECT 0.000 1891.705 18.320 1892.930 ;
        RECT 0.000 1887.870 10.040 1889.095 ;
        RECT 0.000 1887.490 57.880 1887.870 ;
        RECT 0.000 1886.265 1.760 1887.490 ;
        RECT 0.000 1880.825 1.760 1883.655 ;
        RECT 0.000 1875.385 1.760 1878.215 ;
        RECT 0.000 1869.945 1.760 1872.775 ;
        RECT 0.000 1864.505 1.760 1867.335 ;
        RECT 0.000 1859.065 1.760 1861.895 ;
        RECT 0.000 1853.625 1.760 1856.455 ;
        RECT 0.000 1848.185 1.760 1851.015 ;
        RECT 0.000 1842.745 1.760 1845.575 ;
        RECT 0.000 1837.305 1.760 1840.135 ;
        RECT 0.000 1831.865 1.760 1834.695 ;
        RECT 0.000 1826.425 1.760 1829.255 ;
        RECT 0.000 1820.985 1.760 1823.815 ;
        RECT 0.000 1815.545 1.760 1818.375 ;
        RECT 0.000 1810.105 1.760 1812.935 ;
        RECT 0.000 1804.665 1.760 1807.495 ;
        RECT 0.000 1799.225 1.760 1802.055 ;
        RECT 0.000 1793.785 1.760 1796.615 ;
        RECT 0.000 1788.345 1.760 1791.175 ;
        RECT 0.000 1782.905 1.760 1785.735 ;
        RECT 0.000 1777.465 1.760 1780.295 ;
        RECT 0.000 1772.025 1.760 1774.855 ;
        RECT 0.000 1766.585 1.760 1769.415 ;
        RECT 0.000 1761.145 1.760 1763.975 ;
        RECT 0.000 1755.705 1.760 1758.535 ;
        RECT 0.000 1750.265 1.760 1753.095 ;
        RECT 0.000 1744.825 1.760 1747.655 ;
        RECT 0.000 1739.385 1.760 1742.215 ;
        RECT 0.000 1733.945 1.760 1736.775 ;
        RECT 0.000 1728.505 1.760 1731.335 ;
        RECT 0.000 1723.065 1.760 1725.895 ;
        RECT 0.000 1717.625 1.760 1720.455 ;
        RECT 0.000 1712.185 1.760 1715.015 ;
        RECT 0.000 1706.745 1.760 1709.575 ;
        RECT 0.000 1701.305 1.760 1704.135 ;
        RECT 0.000 1695.865 1.760 1698.695 ;
        RECT 0.000 1690.425 1.760 1693.255 ;
        RECT 0.000 1684.985 1.760 1687.815 ;
        RECT 0.000 1679.545 1.760 1682.375 ;
        RECT 0.000 1674.105 1.760 1676.935 ;
        RECT 0.000 1668.665 1.760 1671.495 ;
        RECT 0.000 1663.225 1.760 1666.055 ;
        RECT 0.000 1657.785 1.760 1660.615 ;
        RECT 0.000 1652.345 1.760 1655.175 ;
        RECT 0.000 1646.905 1.760 1649.735 ;
        RECT 0.000 1641.465 1.760 1644.295 ;
        RECT 0.000 1636.025 1.760 1638.855 ;
        RECT 0.000 1630.585 1.760 1633.415 ;
        RECT 0.000 1625.145 1.760 1627.975 ;
        RECT 0.000 1619.705 1.760 1622.535 ;
        RECT 0.000 1614.265 1.760 1617.095 ;
        RECT 0.000 1608.825 1.760 1611.655 ;
        RECT 0.000 1603.385 1.760 1606.215 ;
        RECT 0.000 1597.945 1.760 1600.775 ;
        RECT 0.000 1592.505 1.760 1595.335 ;
        RECT 0.000 1587.065 1.760 1589.895 ;
        RECT 0.000 1581.625 1.760 1584.455 ;
        RECT 0.000 1576.185 1.760 1579.015 ;
        RECT 0.000 1570.745 1.760 1573.575 ;
        RECT 0.000 1565.305 1.760 1568.135 ;
        RECT 0.000 1559.865 1.760 1562.695 ;
        RECT 0.000 1554.425 1.760 1557.255 ;
        RECT 0.000 1548.985 1.760 1551.815 ;
        RECT 0.000 1543.545 1.760 1546.375 ;
        RECT 0.000 1538.105 1.760 1540.935 ;
        RECT 0.000 1532.665 1.760 1535.495 ;
        RECT 0.000 1527.225 1.760 1530.055 ;
        RECT 0.000 1521.785 1.760 1524.615 ;
        RECT 0.000 1516.345 1.760 1519.175 ;
        RECT 0.000 1510.905 1.760 1513.735 ;
        RECT 0.000 1505.465 1.760 1508.295 ;
        RECT 0.000 1500.025 1.760 1502.855 ;
        RECT 0.000 1494.585 1.760 1497.415 ;
        RECT 0.000 1489.145 1.760 1491.975 ;
        RECT 0.000 1483.705 1.760 1486.535 ;
        RECT 0.000 1478.265 1.760 1481.095 ;
        RECT 0.000 1472.825 1.760 1475.655 ;
        RECT 0.000 1467.385 1.760 1470.215 ;
        RECT 0.000 1461.945 1.760 1464.775 ;
        RECT 0.000 1456.505 1.760 1459.335 ;
        RECT 0.000 1451.065 1.760 1453.895 ;
        RECT 0.000 1447.230 14.180 1448.455 ;
        RECT 0.000 1446.850 83.180 1447.230 ;
        RECT 0.000 1445.625 1.760 1446.850 ;
        RECT 0.000 1440.185 1.760 1443.015 ;
        RECT 0.000 1434.745 1.760 1437.575 ;
        RECT 0.000 1429.305 1.760 1432.135 ;
        RECT 0.000 1423.865 1.760 1426.695 ;
        RECT 0.000 1418.425 1.760 1421.255 ;
        RECT 0.000 1412.985 1.760 1415.815 ;
        RECT 0.000 1407.545 1.760 1410.375 ;
        RECT 0.000 1402.105 1.760 1404.935 ;
        RECT 0.000 1396.665 1.760 1399.495 ;
        RECT 0.000 1391.225 1.760 1394.055 ;
        RECT 0.000 1385.785 1.760 1388.615 ;
        RECT 0.000 1380.345 1.760 1383.175 ;
        RECT 0.000 1374.905 1.760 1377.735 ;
        RECT 0.000 1369.465 1.760 1372.295 ;
        RECT 0.000 1364.025 1.760 1366.855 ;
        RECT 0.000 1358.585 1.760 1361.415 ;
        RECT 0.000 1353.145 1.760 1355.975 ;
        RECT 0.000 1347.705 1.760 1350.535 ;
        RECT 0.000 1342.265 1.760 1345.095 ;
        RECT 0.000 1336.825 1.760 1339.655 ;
        RECT 0.000 1331.385 1.760 1334.215 ;
        RECT 0.000 1325.945 1.760 1328.775 ;
        RECT 0.000 1320.505 1.760 1323.335 ;
        RECT 0.000 1315.065 1.760 1317.895 ;
        RECT 0.000 1309.625 1.760 1312.455 ;
        RECT 0.000 1304.185 1.760 1307.015 ;
        RECT 0.000 1298.745 1.760 1301.575 ;
        RECT 0.000 1293.305 1.760 1296.135 ;
        RECT 0.000 1287.865 1.760 1290.695 ;
        RECT 0.000 1282.425 1.760 1285.255 ;
        RECT 0.000 1276.985 1.760 1279.815 ;
        RECT 0.000 1271.545 1.760 1274.375 ;
        RECT 0.000 1266.105 1.760 1268.935 ;
        RECT 0.000 1260.665 1.760 1263.495 ;
        RECT 0.000 1255.225 1.760 1258.055 ;
        RECT 0.000 1249.785 1.760 1252.615 ;
        RECT 0.000 1244.345 1.760 1247.175 ;
        RECT 0.000 1238.905 1.760 1241.735 ;
        RECT 0.000 1233.465 1.760 1236.295 ;
        RECT 0.000 1228.025 1.760 1230.855 ;
        RECT 0.000 1222.585 1.760 1225.415 ;
        RECT 0.000 1217.145 1.760 1219.975 ;
        RECT 0.000 1211.705 1.760 1214.535 ;
        RECT 0.000 1206.265 1.760 1209.095 ;
        RECT 0.000 1200.825 1.760 1203.655 ;
        RECT 0.000 1195.385 1.760 1198.215 ;
        RECT 0.000 1189.945 1.760 1192.775 ;
        RECT 0.000 1184.505 1.760 1187.335 ;
        RECT 0.000 1179.065 1.760 1181.895 ;
        RECT 0.000 1173.625 1.760 1176.455 ;
        RECT 0.000 1168.185 1.760 1171.015 ;
        RECT 0.000 1162.745 1.760 1165.575 ;
        RECT 0.000 1157.305 1.760 1160.135 ;
        RECT 0.000 1151.865 1.760 1154.695 ;
        RECT 0.000 1146.425 1.760 1149.255 ;
        RECT 0.000 1140.985 1.760 1143.815 ;
        RECT 0.000 1135.545 1.760 1138.375 ;
        RECT 0.000 1130.105 1.760 1132.935 ;
        RECT 0.000 1124.665 1.760 1127.495 ;
        RECT 0.000 1119.225 1.760 1122.055 ;
        RECT 0.000 1113.785 1.760 1116.615 ;
        RECT 0.000 1108.345 1.760 1111.175 ;
        RECT 0.000 1102.905 1.760 1105.735 ;
        RECT 0.000 1097.465 1.760 1100.295 ;
        RECT 0.000 1092.025 1.760 1094.855 ;
        RECT 0.000 1086.585 1.760 1089.415 ;
        RECT 0.000 1081.145 1.760 1083.975 ;
        RECT 0.000 1075.705 1.760 1078.535 ;
        RECT 0.000 1070.265 1.760 1073.095 ;
        RECT 0.000 1064.825 1.760 1067.655 ;
        RECT 0.000 1059.385 1.760 1062.215 ;
        RECT 0.000 1053.945 1.760 1056.775 ;
        RECT 0.000 1048.505 1.760 1051.335 ;
        RECT 0.000 1043.065 1.760 1045.895 ;
        RECT 0.000 1037.625 1.760 1040.455 ;
        RECT 0.000 1032.185 1.760 1035.015 ;
        RECT 0.000 1026.745 1.760 1029.575 ;
        RECT 0.000 1021.305 1.760 1024.135 ;
        RECT 0.000 1015.865 1.760 1018.695 ;
        RECT 0.000 1010.425 1.760 1013.255 ;
        RECT 0.000 1004.985 1.760 1007.815 ;
        RECT 0.000 999.545 1.760 1002.375 ;
        RECT 0.000 994.105 1.760 996.935 ;
        RECT 0.000 988.665 1.760 991.495 ;
        RECT 0.000 983.225 1.760 986.055 ;
        RECT 0.000 977.785 1.760 980.615 ;
        RECT 0.000 972.345 1.760 975.175 ;
        RECT 0.000 966.905 1.760 969.735 ;
        RECT 0.000 961.465 1.760 964.295 ;
        RECT 0.000 956.025 1.760 958.855 ;
        RECT 0.000 950.585 1.760 953.415 ;
        RECT 0.000 945.145 1.760 947.975 ;
        RECT 0.000 939.705 1.760 942.535 ;
        RECT 0.000 934.265 1.760 937.095 ;
        RECT 0.000 928.825 1.760 931.655 ;
        RECT 0.000 923.385 1.760 926.215 ;
        RECT 0.000 917.945 1.760 920.775 ;
        RECT 0.000 912.505 1.760 915.335 ;
        RECT 0.000 907.065 1.760 909.895 ;
        RECT 0.000 903.230 1.760 904.455 ;
        RECT 0.000 901.625 10.960 903.230 ;
        RECT 0.000 897.790 9.120 899.015 ;
        RECT 0.000 897.410 15.560 897.790 ;
        RECT 0.000 896.185 1.760 897.410 ;
        RECT 0.000 892.350 9.120 893.575 ;
        RECT 0.000 891.970 28.900 892.350 ;
        RECT 0.000 890.745 1.760 891.970 ;
        RECT 0.000 886.910 14.180 888.135 ;
        RECT 0.000 886.530 16.480 886.910 ;
        RECT 0.000 885.305 1.760 886.530 ;
        RECT 0.000 879.865 1.760 882.695 ;
        RECT 0.000 876.030 1.760 877.255 ;
        RECT 0.000 875.650 41.320 876.030 ;
        RECT 0.000 874.475 9.120 875.650 ;
        RECT 0.000 874.425 2.565 874.475 ;
        RECT 0.000 870.590 1.760 871.815 ;
        RECT 0.000 870.210 26.140 870.590 ;
        RECT 0.000 868.985 13.260 870.210 ;
        RECT 0.000 863.545 1.760 866.375 ;
        RECT 0.000 859.710 1.760 860.935 ;
        RECT 0.000 859.330 75.360 859.710 ;
        RECT 0.000 858.155 9.120 859.330 ;
        RECT 0.000 858.105 2.565 858.155 ;
        RECT 0.000 854.270 1.760 855.495 ;
        RECT 0.000 853.890 167.820 854.270 ;
        RECT 0.000 852.665 20.620 853.890 ;
        RECT 0.000 847.225 1.760 850.055 ;
        RECT 0.000 841.785 1.760 844.615 ;
        RECT 0.000 836.345 1.760 839.175 ;
        RECT 0.000 832.510 1.760 833.735 ;
        RECT 0.000 832.130 123.200 832.510 ;
        RECT 0.000 830.955 18.780 832.130 ;
        RECT 0.000 830.905 2.565 830.955 ;
        RECT 0.000 827.070 1.760 828.295 ;
        RECT 0.000 826.690 19.240 827.070 ;
        RECT 0.000 825.465 17.400 826.690 ;
        RECT 0.000 820.025 1.760 822.855 ;
        RECT 0.000 817.365 2.565 817.415 ;
        RECT 0.000 816.190 9.120 817.365 ;
        RECT 0.000 815.810 19.240 816.190 ;
        RECT 0.000 814.585 1.760 815.810 ;
        RECT 0.000 809.145 1.760 811.975 ;
        RECT 0.000 805.310 1.760 806.535 ;
        RECT 0.000 803.705 10.040 805.310 ;
        RECT 0.000 799.870 14.180 801.095 ;
        RECT 0.000 799.490 15.100 799.870 ;
        RECT 0.000 798.265 1.760 799.490 ;
        RECT 0.000 792.825 1.760 795.655 ;
        RECT 0.000 787.385 1.760 790.215 ;
        RECT 0.000 783.550 9.120 784.775 ;
        RECT 0.000 783.170 84.100 783.550 ;
        RECT 0.000 781.995 10.040 783.170 ;
        RECT 0.000 781.945 2.565 781.995 ;
        RECT 0.000 776.505 1.760 779.335 ;
        RECT 0.000 771.065 1.760 773.895 ;
        RECT 0.000 765.625 1.760 768.455 ;
        RECT 0.000 760.185 1.760 763.015 ;
        RECT 0.000 756.350 1.760 757.575 ;
        RECT 0.000 755.970 476.940 756.350 ;
        RECT 0.000 754.795 27.980 755.970 ;
        RECT 0.000 754.745 2.565 754.795 ;
        RECT 0.000 749.355 10.040 752.135 ;
        RECT 0.000 749.305 2.565 749.355 ;
        RECT 0.000 743.865 1.760 746.695 ;
        RECT 0.000 738.425 16.020 741.255 ;
        RECT 0.000 734.590 13.260 735.815 ;
        RECT 0.000 734.210 268.100 734.590 ;
        RECT 0.000 732.985 1.760 734.210 ;
        RECT 0.000 729.150 1.760 730.375 ;
        RECT 0.000 728.770 19.240 729.150 ;
        RECT 0.000 727.545 18.320 728.770 ;
        RECT 0.000 723.710 1.760 724.935 ;
        RECT 0.000 723.330 178.400 723.710 ;
        RECT 0.000 722.105 27.980 723.330 ;
        RECT 0.000 718.270 1.760 719.495 ;
        RECT 0.000 717.890 180.700 718.270 ;
        RECT 0.000 716.715 41.320 717.890 ;
        RECT 0.000 716.665 2.565 716.715 ;
        RECT 0.000 712.830 1.760 714.055 ;
        RECT 0.000 712.450 237.280 712.830 ;
        RECT 0.000 711.275 9.120 712.450 ;
        RECT 0.000 711.225 2.565 711.275 ;
        RECT 0.000 705.785 1.760 708.615 ;
        RECT 0.000 700.345 1.760 703.175 ;
        RECT 0.000 694.905 1.760 697.735 ;
        RECT 0.000 691.070 14.180 692.295 ;
        RECT 0.000 690.690 72.600 691.070 ;
        RECT 0.000 689.465 17.400 690.690 ;
        RECT 0.000 685.630 1.760 686.855 ;
        RECT 0.000 685.250 125.500 685.630 ;
        RECT 0.000 684.025 10.040 685.250 ;
        RECT 0.000 680.190 14.180 681.415 ;
        RECT 0.000 679.810 126.420 680.190 ;
        RECT 0.000 678.585 1.760 679.810 ;
        RECT 0.000 674.750 14.180 675.975 ;
        RECT 0.000 674.370 350.900 674.750 ;
        RECT 0.000 673.145 1.760 674.370 ;
        RECT 0.000 669.310 1.760 670.535 ;
        RECT 0.000 668.930 166.900 669.310 ;
        RECT 0.000 667.705 9.120 668.930 ;
        RECT 0.000 663.870 14.180 665.095 ;
        RECT 0.000 663.490 23.840 663.870 ;
        RECT 0.000 662.265 1.760 663.490 ;
        RECT 0.000 658.430 14.180 659.655 ;
        RECT 0.000 656.825 23.840 658.430 ;
        RECT 0.000 652.990 14.180 654.215 ;
        RECT 0.000 652.610 41.780 652.990 ;
        RECT 0.000 651.385 10.960 652.610 ;
        RECT 0.000 647.550 14.180 648.775 ;
        RECT 0.000 647.170 41.320 647.550 ;
        RECT 0.000 645.945 1.760 647.170 ;
        RECT 0.000 642.110 14.180 643.335 ;
        RECT 0.000 641.730 84.100 642.110 ;
        RECT 0.000 640.505 1.760 641.730 ;
        RECT 0.000 636.670 14.180 637.895 ;
        RECT 0.000 636.290 71.220 636.670 ;
        RECT 0.000 635.065 1.760 636.290 ;
        RECT 0.000 631.230 1.760 632.455 ;
        RECT 0.000 630.850 105.260 631.230 ;
        RECT 0.000 629.675 16.480 630.850 ;
        RECT 0.000 629.625 2.565 629.675 ;
        RECT 0.000 624.185 1.760 627.015 ;
        RECT 0.000 618.745 1.760 621.575 ;
        RECT 0.000 614.910 14.180 616.135 ;
        RECT 0.000 614.530 251.080 614.910 ;
        RECT 0.000 613.355 25.680 614.530 ;
        RECT 0.000 613.305 9.925 613.355 ;
        RECT 0.000 609.470 1.760 610.695 ;
        RECT 0.000 607.865 20.620 609.470 ;
        RECT 0.000 602.425 1.760 605.255 ;
        RECT 0.000 596.985 1.760 599.815 ;
        RECT 0.000 591.545 1.760 594.375 ;
        RECT 0.000 586.105 1.760 588.935 ;
        RECT 0.000 580.665 1.760 583.495 ;
        RECT 0.000 575.225 1.760 578.055 ;
        RECT 0.000 569.785 1.760 572.615 ;
        RECT 0.000 564.345 1.760 567.175 ;
        RECT 0.000 558.905 1.760 561.735 ;
        RECT 0.000 553.465 1.760 556.295 ;
        RECT 0.000 548.025 1.760 550.855 ;
        RECT 0.000 542.585 1.760 545.415 ;
        RECT 0.000 537.145 1.760 539.975 ;
        RECT 0.000 531.705 1.760 534.535 ;
        RECT 0.000 526.265 1.760 529.095 ;
        RECT 0.000 520.825 1.760 523.655 ;
        RECT 0.000 515.385 1.760 518.215 ;
        RECT 0.000 509.945 1.760 512.775 ;
        RECT 0.000 504.505 1.760 507.335 ;
        RECT 0.000 499.065 1.760 501.895 ;
        RECT 0.000 493.625 1.760 496.455 ;
        RECT 0.000 488.185 1.760 491.015 ;
        RECT 0.000 482.745 1.760 485.575 ;
        RECT 0.000 477.305 1.760 480.135 ;
        RECT 0.000 471.865 1.760 474.695 ;
        RECT 0.000 466.425 1.760 469.255 ;
        RECT 0.000 460.985 1.760 463.815 ;
        RECT 0.000 455.545 1.760 458.375 ;
        RECT 0.000 450.105 1.760 452.935 ;
        RECT 0.000 444.665 1.760 447.495 ;
        RECT 0.000 439.225 1.760 442.055 ;
        RECT 0.000 433.785 1.760 436.615 ;
        RECT 0.000 428.345 1.760 431.175 ;
        RECT 0.000 422.905 1.760 425.735 ;
        RECT 0.000 417.465 1.760 420.295 ;
        RECT 0.000 412.025 1.760 414.855 ;
        RECT 0.000 406.585 1.760 409.415 ;
        RECT 0.000 401.145 1.760 403.975 ;
        RECT 0.000 395.705 1.760 398.535 ;
        RECT 0.000 390.265 1.760 393.095 ;
        RECT 0.000 384.825 1.760 387.655 ;
        RECT 0.000 379.385 1.760 382.215 ;
        RECT 0.000 373.945 1.760 376.775 ;
        RECT 0.000 368.505 1.760 371.335 ;
        RECT 0.000 363.065 1.760 365.895 ;
        RECT 0.000 357.625 1.760 360.455 ;
        RECT 0.000 352.185 1.760 355.015 ;
        RECT 0.000 346.745 1.760 349.575 ;
        RECT 0.000 341.305 1.760 344.135 ;
        RECT 0.000 335.865 1.760 338.695 ;
        RECT 0.000 330.425 1.760 333.255 ;
        RECT 0.000 324.985 1.760 327.815 ;
        RECT 0.000 319.545 1.760 322.375 ;
        RECT 0.000 314.105 1.760 316.935 ;
        RECT 0.000 308.665 1.760 311.495 ;
        RECT 0.000 303.225 1.760 306.055 ;
        RECT 0.000 297.785 1.760 300.615 ;
        RECT 0.000 292.345 1.760 295.175 ;
        RECT 0.000 286.905 1.760 289.735 ;
        RECT 0.000 281.465 1.760 284.295 ;
        RECT 0.000 276.025 1.760 278.855 ;
        RECT 0.000 270.585 1.760 273.415 ;
        RECT 0.000 265.145 1.760 267.975 ;
        RECT 0.000 259.705 1.760 262.535 ;
        RECT 0.000 254.265 1.760 257.095 ;
        RECT 0.000 248.825 1.760 251.655 ;
        RECT 0.000 243.385 1.760 246.215 ;
        RECT 0.000 237.945 1.760 240.775 ;
        RECT 0.000 232.505 1.760 235.335 ;
        RECT 0.000 227.065 1.760 229.895 ;
        RECT 0.000 221.625 1.760 224.455 ;
        RECT 0.000 216.185 1.760 219.015 ;
        RECT 0.000 210.745 1.760 213.575 ;
        RECT 0.000 205.305 1.760 208.135 ;
        RECT 0.000 199.865 1.760 202.695 ;
        RECT 0.000 194.425 1.760 197.255 ;
        RECT 0.000 188.985 1.760 191.815 ;
        RECT 0.000 183.545 1.760 186.375 ;
        RECT 0.000 178.105 1.760 180.935 ;
        RECT 0.000 172.665 1.760 175.495 ;
        RECT 0.000 167.225 1.760 170.055 ;
        RECT 0.000 161.785 1.760 164.615 ;
        RECT 0.000 156.345 1.760 159.175 ;
        RECT 0.000 150.905 1.760 153.735 ;
        RECT 0.000 145.465 1.760 148.295 ;
        RECT 0.000 140.025 1.760 142.855 ;
        RECT 0.000 134.585 1.760 137.415 ;
        RECT 0.000 129.145 1.760 131.975 ;
        RECT 0.000 123.705 1.760 126.535 ;
        RECT 0.000 118.265 1.760 121.095 ;
        RECT 0.000 112.825 1.760 115.655 ;
        RECT 0.000 107.385 1.760 110.215 ;
        RECT 0.000 101.945 1.760 104.775 ;
        RECT 0.000 96.505 1.760 99.335 ;
        RECT 0.000 91.065 1.760 93.895 ;
        RECT 0.000 85.625 1.760 88.455 ;
        RECT 0.000 80.185 1.760 83.015 ;
        RECT 0.000 74.745 1.760 77.575 ;
        RECT 0.000 69.305 1.760 72.135 ;
        RECT 0.000 63.865 1.760 66.695 ;
        RECT 0.000 58.425 1.760 61.255 ;
        RECT 0.000 52.985 1.760 55.815 ;
        RECT 0.000 47.545 1.760 50.375 ;
        RECT 0.000 42.105 1.760 44.935 ;
        RECT 0.000 36.665 1.760 39.495 ;
        RECT 0.000 31.225 1.760 34.055 ;
        RECT 0.000 25.785 1.760 28.615 ;
        RECT 0.000 20.345 1.760 23.175 ;
        RECT 0.000 14.905 1.760 17.735 ;
        RECT 0.000 10.690 1.760 12.295 ;
      LAYER li1 ;
        RECT 0.190 9.945 2889.765 3087.795 ;
      LAYER met1 ;
        RECT 0.190 4.460 2889.825 3087.840 ;
      LAYER met2 ;
        RECT 1.670 4.280 2888.890 3087.870 ;
        RECT 1.670 4.000 11.500 4.280 ;
        RECT 12.340 4.000 46.000 4.280 ;
        RECT 46.840 4.000 80.960 4.280 ;
        RECT 81.800 4.000 115.920 4.280 ;
        RECT 116.760 4.000 150.880 4.280 ;
        RECT 151.720 4.000 185.840 4.280 ;
        RECT 186.680 4.000 220.800 4.280 ;
        RECT 221.640 4.000 255.760 4.280 ;
        RECT 256.600 4.000 290.720 4.280 ;
        RECT 291.560 4.000 325.680 4.280 ;
        RECT 326.520 4.000 360.640 4.280 ;
        RECT 361.480 4.000 395.600 4.280 ;
        RECT 396.440 4.000 430.560 4.280 ;
        RECT 431.400 4.000 465.520 4.280 ;
        RECT 466.360 4.000 500.480 4.280 ;
        RECT 501.320 4.000 535.440 4.280 ;
        RECT 536.280 4.000 570.400 4.280 ;
        RECT 571.240 4.000 605.360 4.280 ;
        RECT 606.200 4.000 640.320 4.280 ;
        RECT 641.160 4.000 675.280 4.280 ;
        RECT 676.120 4.000 710.240 4.280 ;
        RECT 711.080 4.000 744.740 4.280 ;
        RECT 745.580 4.000 779.700 4.280 ;
        RECT 780.540 4.000 814.660 4.280 ;
        RECT 815.500 4.000 849.620 4.280 ;
        RECT 850.460 4.000 884.580 4.280 ;
        RECT 885.420 4.000 919.540 4.280 ;
        RECT 920.380 4.000 954.500 4.280 ;
        RECT 955.340 4.000 989.460 4.280 ;
        RECT 990.300 4.000 1024.420 4.280 ;
        RECT 1025.260 4.000 1059.380 4.280 ;
        RECT 1060.220 4.000 1094.340 4.280 ;
        RECT 1095.180 4.000 1129.300 4.280 ;
        RECT 1130.140 4.000 1164.260 4.280 ;
        RECT 1165.100 4.000 1199.220 4.280 ;
        RECT 1200.060 4.000 1234.180 4.280 ;
        RECT 1235.020 4.000 1269.140 4.280 ;
        RECT 1269.980 4.000 1304.100 4.280 ;
        RECT 1304.940 4.000 1339.060 4.280 ;
        RECT 1339.900 4.000 1374.020 4.280 ;
        RECT 1374.860 4.000 1408.980 4.280 ;
        RECT 1409.820 4.000 1443.940 4.280 ;
        RECT 1444.780 4.000 1478.440 4.280 ;
        RECT 1479.280 4.000 1513.400 4.280 ;
        RECT 1514.240 4.000 1548.360 4.280 ;
        RECT 1549.200 4.000 1583.320 4.280 ;
        RECT 1584.160 4.000 1618.280 4.280 ;
        RECT 1619.120 4.000 1653.240 4.280 ;
        RECT 1654.080 4.000 1688.200 4.280 ;
        RECT 1689.040 4.000 1723.160 4.280 ;
        RECT 1724.000 4.000 1758.120 4.280 ;
        RECT 1758.960 4.000 1793.080 4.280 ;
        RECT 1793.920 4.000 1828.040 4.280 ;
        RECT 1828.880 4.000 1863.000 4.280 ;
        RECT 1863.840 4.000 1897.960 4.280 ;
        RECT 1898.800 4.000 1932.920 4.280 ;
        RECT 1933.760 4.000 1967.880 4.280 ;
        RECT 1968.720 4.000 2002.840 4.280 ;
        RECT 2003.680 4.000 2037.800 4.280 ;
        RECT 2038.640 4.000 2072.760 4.280 ;
        RECT 2073.600 4.000 2107.720 4.280 ;
        RECT 2108.560 4.000 2142.680 4.280 ;
        RECT 2143.520 4.000 2177.640 4.280 ;
        RECT 2178.480 4.000 2212.140 4.280 ;
        RECT 2212.980 4.000 2247.100 4.280 ;
        RECT 2247.940 4.000 2282.060 4.280 ;
        RECT 2282.900 4.000 2317.020 4.280 ;
        RECT 2317.860 4.000 2351.980 4.280 ;
        RECT 2352.820 4.000 2386.940 4.280 ;
        RECT 2387.780 4.000 2421.900 4.280 ;
        RECT 2422.740 4.000 2456.860 4.280 ;
        RECT 2457.700 4.000 2491.820 4.280 ;
        RECT 2492.660 4.000 2526.780 4.280 ;
        RECT 2527.620 4.000 2561.740 4.280 ;
        RECT 2562.580 4.000 2596.700 4.280 ;
        RECT 2597.540 4.000 2631.660 4.280 ;
        RECT 2632.500 4.000 2666.620 4.280 ;
        RECT 2667.460 4.000 2701.580 4.280 ;
        RECT 2702.420 4.000 2736.540 4.280 ;
        RECT 2737.380 4.000 2771.500 4.280 ;
        RECT 2772.340 4.000 2806.460 4.280 ;
        RECT 2807.300 4.000 2841.420 4.280 ;
        RECT 2842.260 4.000 2876.380 4.280 ;
        RECT 2877.220 4.000 2888.890 4.280 ;
      LAYER met3 ;
        RECT 2.555 4.255 2888.005 3087.365 ;
      LAYER met4 ;
        RECT 12.445 10.240 15.310 3082.945 ;
        RECT 17.710 10.240 92.110 3082.945 ;
        RECT 94.510 10.240 168.910 3082.945 ;
        RECT 171.310 10.240 245.710 3082.945 ;
        RECT 248.110 10.240 322.510 3082.945 ;
        RECT 324.910 10.240 399.310 3082.945 ;
        RECT 401.710 10.240 476.110 3082.945 ;
        RECT 478.510 10.240 552.910 3082.945 ;
        RECT 555.310 10.240 629.710 3082.945 ;
        RECT 632.110 10.240 706.510 3082.945 ;
        RECT 708.910 10.240 783.310 3082.945 ;
        RECT 785.710 10.240 860.110 3082.945 ;
        RECT 862.510 10.240 936.910 3082.945 ;
        RECT 939.310 10.240 1013.710 3082.945 ;
        RECT 1016.110 10.240 1090.510 3082.945 ;
        RECT 1092.910 10.240 1167.310 3082.945 ;
        RECT 1169.710 10.240 1244.110 3082.945 ;
        RECT 1246.510 10.240 1320.910 3082.945 ;
        RECT 1323.310 10.240 1397.710 3082.945 ;
        RECT 1400.110 10.240 1474.510 3082.945 ;
        RECT 1476.910 10.240 1551.310 3082.945 ;
        RECT 1553.710 10.240 1628.110 3082.945 ;
        RECT 1630.510 10.240 1704.910 3082.945 ;
        RECT 1707.310 10.240 1781.710 3082.945 ;
        RECT 1784.110 10.240 1858.510 3082.945 ;
        RECT 1860.910 10.240 1935.310 3082.945 ;
        RECT 1937.710 10.240 2012.110 3082.945 ;
        RECT 2014.510 10.240 2088.910 3082.945 ;
        RECT 2091.310 10.240 2165.710 3082.945 ;
        RECT 2168.110 10.240 2242.510 3082.945 ;
        RECT 2244.910 10.240 2319.310 3082.945 ;
        RECT 2321.710 10.240 2396.110 3082.945 ;
        RECT 2398.510 10.240 2472.910 3082.945 ;
        RECT 2475.310 10.240 2549.710 3082.945 ;
        RECT 2552.110 10.240 2626.510 3082.945 ;
        RECT 2628.910 10.240 2703.310 3082.945 ;
        RECT 2705.710 10.240 2780.110 3082.945 ;
        RECT 2782.510 10.240 2856.910 3082.945 ;
        RECT 2859.310 10.240 2875.815 3082.945 ;
        RECT 12.445 9.695 2875.815 10.240 ;
  END
END RAM_6Kx32
END LIBRARY

