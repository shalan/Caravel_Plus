VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM_6Kx32
  CLASS BLOCK ;
  FOREIGN RAM_6Kx32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2889.825 BY 3087.440 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.380 0.000 2247.660 4.000 ;
    END
  END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2596.980 0.000 2597.260 4.000 ;
    END
  END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2631.940 0.000 2632.220 4.000 ;
    END
  END A[11]
  PIN A[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2666.900 0.000 2667.180 4.000 ;
    END
  END A[12]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.340 0.000 2282.620 4.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2317.300 0.000 2317.580 4.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2352.260 0.000 2352.540 4.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2387.220 0.000 2387.500 4.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.180 0.000 2422.460 4.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2457.140 0.000 2457.420 4.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2492.100 0.000 2492.380 4.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.060 0.000 2527.340 4.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.020 0.000 2562.300 4.000 ;
    END
  END A[9]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2701.860 0.000 2702.140 4.000 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.580 0.000 1129.860 4.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.720 0.000 1479.000 4.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.680 0.000 1513.960 4.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.640 0.000 1548.920 4.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.600 0.000 1583.880 4.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.560 0.000 1618.840 4.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.520 0.000 1653.800 4.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.480 0.000 1688.760 4.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.440 0.000 1723.720 4.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.400 0.000 1758.680 4.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.360 0.000 1793.640 4.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.540 0.000 1164.820 4.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.320 0.000 1828.600 4.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.280 0.000 1863.560 4.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.240 0.000 1898.520 4.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.200 0.000 1933.480 4.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1968.160 0.000 1968.440 4.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.120 0.000 2003.400 4.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.080 0.000 2038.360 4.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.040 0.000 2073.320 4.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.000 0.000 2108.280 4.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.960 0.000 2143.240 4.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.500 0.000 1199.780 4.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.920 0.000 2178.200 4.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.420 0.000 2212.700 4.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.460 0.000 1234.740 4.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.420 0.000 1269.700 4.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.380 0.000 1304.660 4.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.340 0.000 1339.620 4.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.300 0.000 1374.580 4.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.260 0.000 1409.540 4.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.220 0.000 1444.500 4.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.780 0.000 12.060 4.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.920 0.000 361.200 4.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.880 0.000 396.160 4.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.840 0.000 431.120 4.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.800 0.000 466.080 4.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.760 0.000 501.040 4.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.720 0.000 536.000 4.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.680 0.000 570.960 4.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.640 0.000 605.920 4.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.600 0.000 640.880 4.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.560 0.000 675.840 4.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.280 0.000 46.560 4.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.520 0.000 710.800 4.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.020 0.000 745.300 4.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.980 0.000 780.260 4.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.940 0.000 815.220 4.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.900 0.000 850.180 4.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.860 0.000 885.140 4.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.820 0.000 920.100 4.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.780 0.000 955.060 4.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.740 0.000 990.020 4.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.700 0.000 1024.980 4.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.240 0.000 81.520 4.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.660 0.000 1059.940 4.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.620 0.000 1094.900 4.000 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.200 0.000 116.480 4.000 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.160 0.000 151.440 4.000 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.120 0.000 186.400 4.000 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.080 0.000 221.360 4.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.040 0.000 256.320 4.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.000 0.000 291.280 4.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.960 0.000 326.240 4.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2876.660 0.000 2876.940 4.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2736.820 0.000 2737.100 4.000 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2771.780 0.000 2772.060 4.000 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2806.740 0.000 2807.020 4.000 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2841.700 0.000 2841.980 4.000 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2780.510 10.640 2782.110 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2626.910 10.640 2628.510 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2473.310 10.640 2474.910 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2319.710 10.640 2321.310 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2166.110 10.640 2167.710 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2012.510 10.640 2014.110 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1858.910 10.640 1860.510 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1705.310 10.640 1706.910 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1551.710 10.640 1553.310 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1398.110 10.640 1399.710 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1244.510 10.640 1246.110 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1090.910 10.640 1092.510 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 937.310 10.640 938.910 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 783.710 10.640 785.310 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 630.110 10.640 631.710 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 476.510 10.640 478.110 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 322.910 10.640 324.510 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 169.310 10.640 170.910 3087.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.710 10.640 17.310 3087.440 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2857.310 10.640 2858.910 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2703.710 10.640 2705.310 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2550.110 10.640 2551.710 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2396.510 10.640 2398.110 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2242.910 10.640 2244.510 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2089.310 10.640 2090.910 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1935.710 10.640 1937.310 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1782.110 10.640 1783.710 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1628.510 10.640 1630.110 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1474.910 10.640 1476.510 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1321.310 10.640 1322.910 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1167.710 10.640 1169.310 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1014.110 10.640 1015.710 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 860.510 10.640 862.110 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 706.910 10.640 708.510 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 553.310 10.640 554.910 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 399.710 10.640 401.310 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.110 10.640 247.710 3087.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 92.510 10.640 94.110 3087.440 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.000 3083.065 2889.180 3085.895 ;
        RECT 0.000 3077.625 2889.180 3080.455 ;
        RECT 0.000 3074.965 1615.325 3075.015 ;
        RECT 0.000 3072.235 2889.180 3074.965 ;
        RECT 0.000 3072.185 1452.485 3072.235 ;
        RECT 0.000 3069.525 904.165 3069.575 ;
        RECT 0.000 3066.795 2889.180 3069.525 ;
        RECT 0.000 3066.745 600.105 3066.795 ;
        RECT 0.000 3064.085 731.205 3064.135 ;
        RECT 0.000 3061.355 2889.180 3064.085 ;
        RECT 0.000 3061.305 555.485 3061.355 ;
        RECT 0.000 3058.645 570.205 3058.695 ;
        RECT 0.000 3055.915 2889.180 3058.645 ;
        RECT 0.000 3055.865 630.465 3055.915 ;
        RECT 0.000 3053.205 773.525 3053.255 ;
        RECT 0.000 3050.475 2889.180 3053.205 ;
        RECT 0.000 3050.425 552.725 3050.475 ;
        RECT 0.000 3047.765 647.025 3047.815 ;
        RECT 0.000 3045.035 2889.180 3047.765 ;
        RECT 0.000 3044.985 667.265 3045.035 ;
        RECT 0.000 3042.325 588.145 3042.375 ;
        RECT 0.000 3039.595 2889.180 3042.325 ;
        RECT 0.000 3039.545 632.765 3039.595 ;
        RECT 0.000 3036.885 569.285 3036.935 ;
        RECT 0.000 3034.155 2889.180 3036.885 ;
        RECT 0.000 3034.105 602.865 3034.155 ;
        RECT 0.000 3031.445 618.045 3031.495 ;
        RECT 0.000 3028.715 2889.180 3031.445 ;
        RECT 0.000 3028.665 562.845 3028.715 ;
        RECT 0.000 3026.005 369.645 3026.055 ;
        RECT 0.000 3023.275 2889.180 3026.005 ;
        RECT 0.000 3023.225 319.505 3023.275 ;
        RECT 0.000 3020.565 278.105 3020.615 ;
        RECT 0.000 3017.835 2889.180 3020.565 ;
        RECT 0.000 3017.785 162.185 3017.835 ;
        RECT 0.000 3015.125 117.565 3015.175 ;
        RECT 0.000 3012.395 2889.180 3015.125 ;
        RECT 0.000 3012.345 99.625 3012.395 ;
        RECT 0.000 3009.685 37.065 3009.735 ;
        RECT 0.000 3006.955 2889.180 3009.685 ;
        RECT 0.000 3006.905 69.725 3006.955 ;
        RECT 0.000 3004.245 55.925 3004.295 ;
        RECT 0.000 3001.515 2889.180 3004.245 ;
        RECT 0.000 3001.465 407.825 3001.515 ;
        RECT 0.000 2998.805 29.245 2998.855 ;
        RECT 0.000 2996.075 2889.180 2998.805 ;
        RECT 0.000 2996.025 11.765 2996.075 ;
        RECT 0.000 2993.365 30.165 2993.415 ;
        RECT 0.000 2990.635 2889.180 2993.365 ;
        RECT 0.000 2990.585 113.885 2990.635 ;
        RECT 0.000 2987.925 57.765 2987.975 ;
        RECT 0.000 2985.195 2889.180 2987.925 ;
        RECT 0.000 2985.145 171.385 2985.195 ;
        RECT 0.000 2982.485 271.205 2982.535 ;
        RECT 0.000 2979.755 2889.180 2982.485 ;
        RECT 0.000 2979.705 3.485 2979.755 ;
        RECT 0.000 2977.045 36.605 2977.095 ;
        RECT 0.000 2974.315 2889.180 2977.045 ;
        RECT 0.000 2974.265 98.245 2974.315 ;
        RECT 0.000 2971.605 147.925 2971.655 ;
        RECT 0.000 2968.875 2889.180 2971.605 ;
        RECT 0.000 2968.825 283.625 2968.875 ;
        RECT 0.000 2966.165 8.545 2966.215 ;
        RECT 0.000 2963.435 2889.180 2966.165 ;
        RECT 0.000 2963.385 67.885 2963.435 ;
        RECT 0.000 2960.725 380.685 2960.775 ;
        RECT 0.000 2957.995 2889.180 2960.725 ;
        RECT 0.000 2957.945 2.565 2957.995 ;
        RECT 0.000 2955.285 117.105 2955.335 ;
        RECT 0.000 2952.555 2889.180 2955.285 ;
        RECT 0.000 2952.505 43.505 2952.555 ;
        RECT 0.000 2949.845 224.285 2949.895 ;
        RECT 0.000 2947.115 2889.180 2949.845 ;
        RECT 0.000 2947.065 115.725 2947.115 ;
        RECT 0.000 2944.405 100.085 2944.455 ;
        RECT 0.000 2941.675 2889.180 2944.405 ;
        RECT 0.000 2941.625 31.545 2941.675 ;
        RECT 0.000 2938.965 72.485 2939.015 ;
        RECT 0.000 2936.235 2889.180 2938.965 ;
        RECT 0.000 2936.185 154.365 2936.235 ;
        RECT 0.000 2933.525 2.565 2933.575 ;
        RECT 0.000 2930.795 2889.180 2933.525 ;
        RECT 0.000 2930.745 87.205 2930.795 ;
        RECT 0.000 2928.085 273.045 2928.135 ;
        RECT 0.000 2925.355 2889.180 2928.085 ;
        RECT 0.000 2925.305 3.945 2925.355 ;
        RECT 0.000 2922.645 52.245 2922.695 ;
        RECT 0.000 2919.915 2889.180 2922.645 ;
        RECT 0.000 2919.865 219.225 2919.915 ;
        RECT 0.000 2917.205 34.765 2917.255 ;
        RECT 0.000 2914.475 2889.180 2917.205 ;
        RECT 0.000 2914.425 68.345 2914.475 ;
        RECT 0.000 2911.765 110.665 2911.815 ;
        RECT 0.000 2909.035 2889.180 2911.765 ;
        RECT 0.000 2908.985 20.965 2909.035 ;
        RECT 0.000 2906.325 279.485 2906.375 ;
        RECT 0.000 2903.595 2889.180 2906.325 ;
        RECT 0.000 2903.545 236.245 2903.595 ;
        RECT 0.000 2900.885 24.645 2900.935 ;
        RECT 0.000 2898.155 2889.180 2900.885 ;
        RECT 0.000 2898.105 96.405 2898.155 ;
        RECT 0.000 2895.445 9.005 2895.495 ;
        RECT 0.000 2892.715 2889.180 2895.445 ;
        RECT 0.000 2892.665 90.425 2892.715 ;
        RECT 0.000 2890.005 303.865 2890.055 ;
        RECT 0.000 2887.275 2889.180 2890.005 ;
        RECT 0.000 2887.225 21.425 2887.275 ;
        RECT 0.000 2884.565 205.425 2884.615 ;
        RECT 0.000 2881.835 2889.180 2884.565 ;
        RECT 0.000 2881.785 71.105 2881.835 ;
        RECT 0.000 2879.125 131.365 2879.175 ;
        RECT 0.000 2876.395 2889.180 2879.125 ;
        RECT 0.000 2876.345 38.905 2876.395 ;
        RECT 0.000 2873.685 6.245 2873.735 ;
        RECT 0.000 2870.955 2889.180 2873.685 ;
        RECT 0.000 2870.905 486.485 2870.955 ;
        RECT 0.000 2868.245 278.105 2868.295 ;
        RECT 0.000 2865.515 2889.180 2868.245 ;
        RECT 0.000 2865.465 296.505 2865.515 ;
        RECT 0.000 2862.805 233.485 2862.855 ;
        RECT 0.000 2860.075 2889.180 2862.805 ;
        RECT 0.000 2860.025 3.945 2860.075 ;
        RECT 0.000 2857.365 79.385 2857.415 ;
        RECT 0.000 2854.635 2889.180 2857.365 ;
        RECT 0.000 2854.585 423.465 2854.635 ;
        RECT 0.000 2851.925 72.025 2851.975 ;
        RECT 0.000 2849.195 2889.180 2851.925 ;
        RECT 0.000 2849.145 9.925 2849.195 ;
        RECT 0.000 2846.485 37.065 2846.535 ;
        RECT 0.000 2843.755 2889.180 2846.485 ;
        RECT 0.000 2843.705 21.425 2843.755 ;
        RECT 0.000 2841.045 54.545 2841.095 ;
        RECT 0.000 2838.315 2889.180 2841.045 ;
        RECT 0.000 2838.265 37.525 2838.315 ;
        RECT 0.000 2835.605 302.485 2835.655 ;
        RECT 0.000 2832.875 2889.180 2835.605 ;
        RECT 0.000 2832.825 129.065 2832.875 ;
        RECT 0.000 2830.165 2.565 2830.215 ;
        RECT 0.000 2827.435 2889.180 2830.165 ;
        RECT 0.000 2827.385 77.085 2827.435 ;
        RECT 0.000 2824.725 90.425 2824.775 ;
        RECT 0.000 2821.995 2889.180 2824.725 ;
        RECT 0.000 2821.945 246.365 2821.995 ;
        RECT 0.000 2819.285 9.005 2819.335 ;
        RECT 0.000 2816.555 2889.180 2819.285 ;
        RECT 0.000 2816.505 106.985 2816.555 ;
        RECT 0.000 2813.845 129.065 2813.895 ;
        RECT 0.000 2811.115 2889.180 2813.845 ;
        RECT 0.000 2811.065 114.805 2811.115 ;
        RECT 0.000 2808.405 55.465 2808.455 ;
        RECT 0.000 2805.675 2889.180 2808.405 ;
        RECT 0.000 2805.625 59.145 2805.675 ;
        RECT 0.000 2802.965 20.505 2803.015 ;
        RECT 0.000 2800.235 2889.180 2802.965 ;
        RECT 0.000 2800.185 102.845 2800.235 ;
        RECT 0.000 2797.525 7.165 2797.575 ;
        RECT 0.000 2794.795 2889.180 2797.525 ;
        RECT 0.000 2794.745 177.825 2794.795 ;
        RECT 0.000 2792.085 23.265 2792.135 ;
        RECT 0.000 2789.355 2889.180 2792.085 ;
        RECT 0.000 2789.305 66.965 2789.355 ;
        RECT 0.000 2786.645 51.785 2786.695 ;
        RECT 0.000 2783.915 2889.180 2786.645 ;
        RECT 0.000 2783.865 106.985 2783.915 ;
        RECT 0.000 2781.205 3.945 2781.255 ;
        RECT 0.000 2778.475 2889.180 2781.205 ;
        RECT 0.000 2778.425 37.525 2778.475 ;
        RECT 0.000 2775.765 177.365 2775.815 ;
        RECT 0.000 2773.035 2889.180 2775.765 ;
        RECT 0.000 2772.985 275.345 2773.035 ;
        RECT 0.000 2770.325 115.725 2770.375 ;
        RECT 0.000 2767.595 2889.180 2770.325 ;
        RECT 0.000 2767.545 327.785 2767.595 ;
        RECT 0.000 2764.885 8.085 2764.935 ;
        RECT 0.000 2762.155 2889.180 2764.885 ;
        RECT 0.000 2762.105 22.805 2762.155 ;
        RECT 0.000 2759.445 363.205 2759.495 ;
        RECT 0.000 2756.715 2889.180 2759.445 ;
        RECT 0.000 2756.665 77.085 2756.715 ;
        RECT 0.000 2754.005 105.605 2754.055 ;
        RECT 0.000 2751.275 2889.180 2754.005 ;
        RECT 0.000 2751.225 22.805 2751.275 ;
        RECT 0.000 2748.565 132.285 2748.615 ;
        RECT 0.000 2745.835 2889.180 2748.565 ;
        RECT 0.000 2745.785 40.285 2745.835 ;
        RECT 0.000 2743.125 37.065 2743.175 ;
        RECT 0.000 2740.395 2889.180 2743.125 ;
        RECT 0.000 2740.345 4.865 2740.395 ;
        RECT 0.000 2737.685 187.485 2737.735 ;
        RECT 0.000 2734.955 2889.180 2737.685 ;
        RECT 0.000 2734.905 89.045 2734.955 ;
        RECT 0.000 2732.245 27.405 2732.295 ;
        RECT 0.000 2729.515 2889.180 2732.245 ;
        RECT 0.000 2729.465 115.265 2729.515 ;
        RECT 0.000 2726.805 20.505 2726.855 ;
        RECT 0.000 2724.075 2889.180 2726.805 ;
        RECT 0.000 2724.025 103.765 2724.075 ;
        RECT 0.000 2721.365 43.965 2721.415 ;
        RECT 0.000 2718.635 2889.180 2721.365 ;
        RECT 0.000 2718.585 153.905 2718.635 ;
        RECT 0.000 2715.925 213.245 2715.975 ;
        RECT 0.000 2713.195 2889.180 2715.925 ;
        RECT 0.000 2713.145 405.525 2713.195 ;
        RECT 0.000 2710.485 56.385 2710.535 ;
        RECT 0.000 2707.755 2889.180 2710.485 ;
        RECT 0.000 2707.705 163.105 2707.755 ;
        RECT 0.000 2705.045 26.025 2705.095 ;
        RECT 0.000 2702.315 2889.180 2705.045 ;
        RECT 0.000 2702.265 93.185 2702.315 ;
        RECT 0.000 2699.605 37.065 2699.655 ;
        RECT 0.000 2696.875 2889.180 2699.605 ;
        RECT 0.000 2696.825 176.905 2696.875 ;
        RECT 0.000 2694.165 9.005 2694.215 ;
        RECT 0.000 2691.435 2889.180 2694.165 ;
        RECT 0.000 2691.385 114.345 2691.435 ;
        RECT 0.000 2688.725 27.865 2688.775 ;
        RECT 0.000 2685.995 2889.180 2688.725 ;
        RECT 0.000 2685.945 76.165 2685.995 ;
        RECT 0.000 2683.285 472.225 2683.335 ;
        RECT 0.000 2680.555 2889.180 2683.285 ;
        RECT 0.000 2680.505 394.485 2680.555 ;
        RECT 0.000 2677.845 326.405 2677.895 ;
        RECT 0.000 2675.115 2889.180 2677.845 ;
        RECT 0.000 2675.065 692.105 2675.115 ;
        RECT 0.000 2672.405 313.525 2672.455 ;
        RECT 0.000 2669.675 2889.180 2672.405 ;
        RECT 0.000 2669.625 359.525 2669.675 ;
        RECT 0.000 2666.965 195.765 2667.015 ;
        RECT 0.000 2664.235 2889.180 2666.965 ;
        RECT 0.000 2664.185 94.565 2664.235 ;
        RECT 0.000 2661.525 26.945 2661.575 ;
        RECT 0.000 2658.795 2889.180 2661.525 ;
        RECT 0.000 2658.745 155.285 2658.795 ;
        RECT 0.000 2656.085 45.805 2656.135 ;
        RECT 0.000 2653.355 2889.180 2656.085 ;
        RECT 0.000 2653.305 129.065 2653.355 ;
        RECT 0.000 2650.645 26.485 2650.695 ;
        RECT 0.000 2647.915 2889.180 2650.645 ;
        RECT 0.000 2647.865 95.945 2647.915 ;
        RECT 0.000 2645.205 26.485 2645.255 ;
        RECT 0.000 2642.475 2889.180 2645.205 ;
        RECT 0.000 2642.425 127.685 2642.475 ;
        RECT 0.000 2639.765 37.065 2639.815 ;
        RECT 0.000 2637.035 2889.180 2639.765 ;
        RECT 0.000 2636.985 57.765 2637.035 ;
        RECT 0.000 2634.325 23.725 2634.375 ;
        RECT 0.000 2631.595 2889.180 2634.325 ;
        RECT 0.000 2631.545 118.485 2631.595 ;
        RECT 0.000 2628.885 218.765 2628.935 ;
        RECT 0.000 2626.155 2889.180 2628.885 ;
        RECT 0.000 2626.105 86.745 2626.155 ;
        RECT 0.000 2623.445 23.265 2623.495 ;
        RECT 0.000 2620.715 2889.180 2623.445 ;
        RECT 0.000 2620.665 127.685 2620.715 ;
        RECT 0.000 2618.005 65.125 2618.055 ;
        RECT 0.000 2615.275 2889.180 2618.005 ;
        RECT 0.000 2615.225 269.825 2615.275 ;
        RECT 0.000 2612.565 36.605 2612.615 ;
        RECT 0.000 2609.835 2889.180 2612.565 ;
        RECT 0.000 2609.785 22.805 2609.835 ;
        RECT 0.000 2607.125 26.025 2607.175 ;
        RECT 0.000 2604.395 2889.180 2607.125 ;
        RECT 0.000 2604.345 290.525 2604.395 ;
        RECT 0.000 2601.685 467.165 2601.735 ;
        RECT 0.000 2598.955 2889.180 2601.685 ;
        RECT 0.000 2598.905 198.065 2598.955 ;
        RECT 0.000 2596.245 56.845 2596.295 ;
        RECT 0.000 2593.515 2889.180 2596.245 ;
        RECT 0.000 2593.465 42.585 2593.515 ;
        RECT 0.000 2590.805 131.825 2590.855 ;
        RECT 0.000 2588.075 2889.180 2590.805 ;
        RECT 0.000 2588.025 29.705 2588.075 ;
        RECT 0.000 2585.365 28.325 2585.415 ;
        RECT 0.000 2582.635 2889.180 2585.365 ;
        RECT 0.000 2582.585 119.865 2582.635 ;
        RECT 0.000 2579.925 230.725 2579.975 ;
        RECT 0.000 2577.195 2889.180 2579.925 ;
        RECT 0.000 2577.145 415.645 2577.195 ;
        RECT 0.000 2574.485 26.485 2574.535 ;
        RECT 0.000 2571.755 2889.180 2574.485 ;
        RECT 0.000 2571.705 442.785 2571.755 ;
        RECT 0.000 2569.045 107.905 2569.095 ;
        RECT 0.000 2566.315 2889.180 2569.045 ;
        RECT 0.000 2566.265 22.805 2566.315 ;
        RECT 0.000 2563.605 141.485 2563.655 ;
        RECT 0.000 2560.875 2889.180 2563.605 ;
        RECT 0.000 2560.825 66.965 2560.875 ;
        RECT 0.000 2558.165 25.565 2558.215 ;
        RECT 0.000 2555.435 2889.180 2558.165 ;
        RECT 0.000 2555.385 43.505 2555.435 ;
        RECT 0.000 2552.725 393.105 2552.775 ;
        RECT 0.000 2549.995 2889.180 2552.725 ;
        RECT 0.000 2549.945 38.445 2549.995 ;
        RECT 0.000 2547.285 56.385 2547.335 ;
        RECT 0.000 2544.555 2889.180 2547.285 ;
        RECT 0.000 2544.505 175.065 2544.555 ;
        RECT 0.000 2541.845 24.645 2541.895 ;
        RECT 0.000 2539.115 2889.180 2541.845 ;
        RECT 0.000 2539.065 219.225 2539.115 ;
        RECT 0.000 2536.405 136.425 2536.455 ;
        RECT 0.000 2533.675 2889.180 2536.405 ;
        RECT 0.000 2533.625 57.765 2533.675 ;
        RECT 0.000 2530.965 23.265 2531.015 ;
        RECT 0.000 2528.235 2889.180 2530.965 ;
        RECT 0.000 2528.185 302.945 2528.235 ;
        RECT 0.000 2525.525 288.225 2525.575 ;
        RECT 0.000 2522.795 2889.180 2525.525 ;
        RECT 0.000 2522.745 22.805 2522.795 ;
        RECT 0.000 2520.085 87.665 2520.135 ;
        RECT 0.000 2517.355 2889.180 2520.085 ;
        RECT 0.000 2517.305 50.865 2517.355 ;
        RECT 0.000 2514.645 105.145 2514.695 ;
        RECT 0.000 2511.915 2889.180 2514.645 ;
        RECT 0.000 2511.865 22.805 2511.915 ;
        RECT 0.000 2509.205 177.365 2509.255 ;
        RECT 0.000 2506.475 2889.180 2509.205 ;
        RECT 0.000 2506.425 434.965 2506.475 ;
        RECT 0.000 2503.765 652.545 2503.815 ;
        RECT 0.000 2501.035 2889.180 2503.765 ;
        RECT 0.000 2500.985 575.265 2501.035 ;
        RECT 0.000 2498.325 1325.065 2498.375 ;
        RECT 0.000 2495.595 2889.180 2498.325 ;
        RECT 0.000 2495.545 50.865 2495.595 ;
        RECT 0.000 2492.885 268.905 2492.935 ;
        RECT 0.000 2490.155 2889.180 2492.885 ;
        RECT 0.000 2490.105 78.925 2490.155 ;
        RECT 0.000 2487.445 4.405 2487.495 ;
        RECT 0.000 2484.715 2889.180 2487.445 ;
        RECT 0.000 2484.665 19.125 2484.715 ;
        RECT 0.000 2482.005 117.565 2482.055 ;
        RECT 0.000 2479.275 2889.180 2482.005 ;
        RECT 0.000 2479.225 71.105 2479.275 ;
        RECT 0.000 2476.565 296.505 2476.615 ;
        RECT 0.000 2473.835 2889.180 2476.565 ;
        RECT 0.000 2473.785 20.505 2473.835 ;
        RECT 0.000 2471.125 84.445 2471.175 ;
        RECT 0.000 2468.395 2889.180 2471.125 ;
        RECT 0.000 2468.345 261.545 2468.395 ;
        RECT 0.000 2465.685 4.405 2465.735 ;
        RECT 0.000 2462.955 2889.180 2465.685 ;
        RECT 0.000 2462.905 37.985 2462.955 ;
        RECT 0.000 2460.245 224.285 2460.295 ;
        RECT 0.000 2457.515 2889.180 2460.245 ;
        RECT 0.000 2457.465 22.805 2457.515 ;
        RECT 0.000 2454.805 184.265 2454.855 ;
        RECT 0.000 2452.075 2889.180 2454.805 ;
        RECT 0.000 2452.025 3.485 2452.075 ;
        RECT 0.000 2449.365 141.025 2449.415 ;
        RECT 0.000 2446.635 2889.180 2449.365 ;
        RECT 0.000 2446.585 37.525 2446.635 ;
        RECT 0.000 2443.925 21.425 2443.975 ;
        RECT 0.000 2441.195 2889.180 2443.925 ;
        RECT 0.000 2441.145 3.945 2441.195 ;
        RECT 0.000 2438.485 88.125 2438.535 ;
        RECT 0.000 2435.755 2889.180 2438.485 ;
        RECT 0.000 2435.705 69.725 2435.755 ;
        RECT 0.000 2433.045 130.445 2433.095 ;
        RECT 0.000 2430.315 2889.180 2433.045 ;
        RECT 0.000 2430.265 160.805 2430.315 ;
        RECT 0.000 2427.605 44.885 2427.655 ;
        RECT 0.000 2424.875 2889.180 2427.605 ;
        RECT 0.000 2424.825 210.945 2424.875 ;
        RECT 0.000 2422.165 3.945 2422.215 ;
        RECT 0.000 2419.435 2889.180 2422.165 ;
        RECT 0.000 2419.385 22.805 2419.435 ;
        RECT 0.000 2416.725 121.245 2416.775 ;
        RECT 0.000 2413.995 2889.180 2416.725 ;
        RECT 0.000 2413.945 341.585 2413.995 ;
        RECT 0.000 2411.285 92.725 2411.335 ;
        RECT 0.000 2408.555 2889.180 2411.285 ;
        RECT 0.000 2408.505 156.205 2408.555 ;
        RECT 0.000 2405.845 420.705 2405.895 ;
        RECT 0.000 2403.115 2889.180 2405.845 ;
        RECT 0.000 2403.065 18.665 2403.115 ;
        RECT 0.000 2400.405 5.325 2400.455 ;
        RECT 0.000 2397.675 2889.180 2400.405 ;
        RECT 0.000 2397.625 121.245 2397.675 ;
        RECT 0.000 2394.965 75.705 2395.015 ;
        RECT 0.000 2392.235 2889.180 2394.965 ;
        RECT 0.000 2392.185 406.905 2392.235 ;
        RECT 0.000 2389.525 61.905 2389.575 ;
        RECT 0.000 2386.795 2889.180 2389.525 ;
        RECT 0.000 2386.745 22.805 2386.795 ;
        RECT 0.000 2384.085 120.785 2384.135 ;
        RECT 0.000 2381.355 2889.180 2384.085 ;
        RECT 0.000 2381.305 42.125 2381.355 ;
        RECT 0.000 2378.645 6.245 2378.695 ;
        RECT 0.000 2375.915 2889.180 2378.645 ;
        RECT 0.000 2375.865 562.845 2375.915 ;
        RECT 0.000 2373.205 61.445 2373.255 ;
        RECT 0.000 2370.475 2889.180 2373.205 ;
        RECT 0.000 2370.425 216.465 2370.475 ;
        RECT 0.000 2367.765 44.425 2367.815 ;
        RECT 0.000 2365.035 2889.180 2367.765 ;
        RECT 0.000 2364.985 10.385 2365.035 ;
        RECT 0.000 2362.325 26.945 2362.375 ;
        RECT 0.000 2359.595 2889.180 2362.325 ;
        RECT 0.000 2359.545 267.525 2359.595 ;
        RECT 0.000 2356.885 89.505 2356.935 ;
        RECT 0.000 2354.155 2889.180 2356.885 ;
        RECT 0.000 2354.105 188.865 2354.155 ;
        RECT 0.000 2351.445 23.265 2351.495 ;
        RECT 0.000 2348.715 2889.180 2351.445 ;
        RECT 0.000 2348.665 40.745 2348.715 ;
        RECT 0.000 2346.005 121.245 2346.055 ;
        RECT 0.000 2343.275 2889.180 2346.005 ;
        RECT 0.000 2343.225 3.485 2343.275 ;
        RECT 0.000 2340.565 93.185 2340.615 ;
        RECT 0.000 2337.835 2889.180 2340.565 ;
        RECT 0.000 2337.785 142.405 2337.835 ;
        RECT 0.000 2335.125 457.505 2335.175 ;
        RECT 0.000 2332.395 2889.180 2335.125 ;
        RECT 0.000 2332.345 161.725 2332.395 ;
        RECT 0.000 2329.685 175.525 2329.735 ;
        RECT 0.000 2326.955 2889.180 2329.685 ;
        RECT 0.000 2326.905 78.925 2326.955 ;
        RECT 0.000 2324.245 3.945 2324.295 ;
        RECT 0.000 2321.515 2889.180 2324.245 ;
        RECT 0.000 2321.465 19.125 2321.515 ;
        RECT 0.000 2318.805 53.165 2318.855 ;
        RECT 0.000 2316.075 2889.180 2318.805 ;
        RECT 0.000 2316.025 37.985 2316.075 ;
        RECT 0.000 2313.365 8.545 2313.415 ;
        RECT 0.000 2310.635 2889.180 2313.365 ;
        RECT 0.000 2310.585 338.365 2310.635 ;
        RECT 0.000 2307.925 501.205 2307.975 ;
        RECT 0.000 2305.195 2889.180 2307.925 ;
        RECT 0.000 2305.145 443.705 2305.195 ;
        RECT 0.000 2302.485 305.245 2302.535 ;
        RECT 0.000 2299.755 2889.180 2302.485 ;
        RECT 0.000 2299.705 675.085 2299.755 ;
        RECT 0.000 2297.045 84.905 2297.095 ;
        RECT 0.000 2294.315 2889.180 2297.045 ;
        RECT 0.000 2294.265 2.565 2294.315 ;
        RECT 0.000 2291.605 72.025 2291.655 ;
        RECT 0.000 2288.875 2889.180 2291.605 ;
        RECT 0.000 2288.825 43.045 2288.875 ;
        RECT 0.000 2286.165 27.865 2286.215 ;
        RECT 0.000 2283.435 2889.180 2286.165 ;
        RECT 0.000 2283.385 43.965 2283.435 ;
        RECT 0.000 2280.725 149.305 2280.775 ;
        RECT 0.000 2277.995 2889.180 2280.725 ;
        RECT 0.000 2277.945 133.205 2277.995 ;
        RECT 0.000 2275.285 15.905 2275.335 ;
        RECT 0.000 2272.555 2889.180 2275.285 ;
        RECT 0.000 2272.505 116.645 2272.555 ;
        RECT 0.000 2269.845 28.785 2269.895 ;
        RECT 0.000 2267.115 2889.180 2269.845 ;
        RECT 0.000 2267.065 149.765 2267.115 ;
        RECT 0.000 2264.405 74.325 2264.455 ;
        RECT 0.000 2261.675 2889.180 2264.405 ;
        RECT 0.000 2261.625 10.845 2261.675 ;
        RECT 0.000 2258.965 48.105 2259.015 ;
        RECT 0.000 2256.235 2889.180 2258.965 ;
        RECT 0.000 2256.185 135.045 2256.235 ;
        RECT 0.000 2253.525 72.025 2253.575 ;
        RECT 0.000 2250.795 2889.180 2253.525 ;
        RECT 0.000 2250.745 86.285 2250.795 ;
        RECT 0.000 2248.085 289.605 2248.135 ;
        RECT 0.000 2245.355 2889.180 2248.085 ;
        RECT 0.000 2245.305 5.785 2245.355 ;
        RECT 0.000 2242.645 37.065 2242.695 ;
        RECT 0.000 2239.915 2889.180 2242.645 ;
        RECT 0.000 2239.865 22.345 2239.915 ;
        RECT 0.000 2237.205 331.925 2237.255 ;
        RECT 0.000 2234.475 2889.180 2237.205 ;
        RECT 0.000 2234.425 87.205 2234.475 ;
        RECT 0.000 2231.765 6.705 2231.815 ;
        RECT 0.000 2229.035 2889.180 2231.765 ;
        RECT 0.000 2228.985 331.465 2229.035 ;
        RECT 0.000 2226.325 72.485 2226.375 ;
        RECT 0.000 2223.595 2889.180 2226.325 ;
        RECT 0.000 2223.545 39.825 2223.595 ;
        RECT 0.000 2220.885 25.565 2220.935 ;
        RECT 0.000 2218.155 2889.180 2220.885 ;
        RECT 0.000 2218.105 133.205 2218.155 ;
        RECT 0.000 2215.445 101.005 2215.495 ;
        RECT 0.000 2212.715 2889.180 2215.445 ;
        RECT 0.000 2212.665 345.725 2212.715 ;
        RECT 0.000 2210.005 261.085 2210.055 ;
        RECT 0.000 2207.275 2889.180 2210.005 ;
        RECT 0.000 2207.225 3.945 2207.275 ;
        RECT 0.000 2204.565 147.925 2204.615 ;
        RECT 0.000 2201.835 2889.180 2204.565 ;
        RECT 0.000 2201.785 340.205 2201.835 ;
        RECT 0.000 2199.125 54.085 2199.175 ;
        RECT 0.000 2196.395 2889.180 2199.125 ;
        RECT 0.000 2196.345 8.545 2196.395 ;
        RECT 0.000 2193.685 214.625 2193.735 ;
        RECT 0.000 2190.955 2889.180 2193.685 ;
        RECT 0.000 2190.905 22.805 2190.955 ;
        RECT 0.000 2188.245 65.125 2188.295 ;
        RECT 0.000 2185.515 2889.180 2188.245 ;
        RECT 0.000 2185.465 133.665 2185.515 ;
        RECT 0.000 2182.805 276.265 2182.855 ;
        RECT 0.000 2180.075 2889.180 2182.805 ;
        RECT 0.000 2180.025 49.485 2180.075 ;
        RECT 0.000 2177.365 93.185 2177.415 ;
        RECT 0.000 2174.635 2889.180 2177.365 ;
        RECT 0.000 2174.585 4.865 2174.635 ;
        RECT 0.000 2171.925 164.945 2171.975 ;
        RECT 0.000 2169.195 2889.180 2171.925 ;
        RECT 0.000 2169.145 115.265 2169.195 ;
        RECT 0.000 2166.485 75.245 2166.535 ;
        RECT 0.000 2163.755 2889.180 2166.485 ;
        RECT 0.000 2163.705 22.805 2163.755 ;
        RECT 0.000 2161.045 9.005 2161.095 ;
        RECT 0.000 2158.315 2889.180 2161.045 ;
        RECT 0.000 2158.265 241.765 2158.315 ;
        RECT 0.000 2155.605 164.945 2155.655 ;
        RECT 0.000 2152.875 2889.180 2155.605 ;
        RECT 0.000 2152.825 144.705 2152.875 ;
        RECT 0.000 2150.165 43.965 2150.215 ;
        RECT 0.000 2147.435 2889.180 2150.165 ;
        RECT 0.000 2147.385 123.085 2147.435 ;
        RECT 0.000 2144.725 57.765 2144.775 ;
        RECT 0.000 2141.995 2889.180 2144.725 ;
        RECT 0.000 2141.945 21.425 2141.995 ;
        RECT 0.000 2139.285 9.005 2139.335 ;
        RECT 0.000 2136.555 2889.180 2139.285 ;
        RECT 0.000 2136.505 37.065 2136.555 ;
        RECT 0.000 2133.845 612.985 2133.895 ;
        RECT 0.000 2131.115 2889.180 2133.845 ;
        RECT 0.000 2131.065 238.085 2131.115 ;
        RECT 0.000 2128.405 233.485 2128.455 ;
        RECT 0.000 2125.675 2889.180 2128.405 ;
        RECT 0.000 2125.625 376.085 2125.675 ;
        RECT 0.000 2122.965 315.365 2123.015 ;
        RECT 0.000 2120.235 2889.180 2122.965 ;
        RECT 0.000 2120.185 275.345 2120.235 ;
        RECT 0.000 2117.525 249.585 2117.575 ;
        RECT 0.000 2114.795 2889.180 2117.525 ;
        RECT 0.000 2114.745 96.865 2114.795 ;
        RECT 0.000 2112.085 166.785 2112.135 ;
        RECT 0.000 2109.355 2889.180 2112.085 ;
        RECT 0.000 2109.305 78.925 2109.355 ;
        RECT 0.000 2106.645 112.505 2106.695 ;
        RECT 0.000 2103.915 2889.180 2106.645 ;
        RECT 0.000 2103.865 127.685 2103.915 ;
        RECT 0.000 2101.205 144.705 2101.255 ;
        RECT 0.000 2098.475 2889.180 2101.205 ;
        RECT 0.000 2098.425 32.925 2098.475 ;
        RECT 0.000 2095.765 49.485 2095.815 ;
        RECT 0.000 2093.035 2889.180 2095.765 ;
        RECT 0.000 2092.985 233.485 2093.035 ;
        RECT 0.000 2090.325 278.105 2090.375 ;
        RECT 0.000 2087.595 2889.180 2090.325 ;
        RECT 0.000 2087.545 5.325 2087.595 ;
        RECT 0.000 2084.885 44.885 2084.935 ;
        RECT 0.000 2082.155 2889.180 2084.885 ;
        RECT 0.000 2082.105 170.005 2082.155 ;
        RECT 0.000 2079.445 61.905 2079.495 ;
        RECT 0.000 2076.715 2889.180 2079.445 ;
        RECT 0.000 2076.665 97.785 2076.715 ;
        RECT 0.000 2074.005 338.365 2074.055 ;
        RECT 0.000 2071.275 2889.180 2074.005 ;
        RECT 0.000 2071.225 413.805 2071.275 ;
        RECT 0.000 2068.565 80.765 2068.615 ;
        RECT 0.000 2065.835 2889.180 2068.565 ;
        RECT 0.000 2065.785 4.405 2065.835 ;
        RECT 0.000 2063.125 29.705 2063.175 ;
        RECT 0.000 2060.395 2889.180 2063.125 ;
        RECT 0.000 2060.345 125.385 2060.395 ;
        RECT 0.000 2057.685 49.485 2057.735 ;
        RECT 0.000 2054.955 2889.180 2057.685 ;
        RECT 0.000 2054.905 62.825 2054.955 ;
        RECT 0.000 2052.245 363.665 2052.295 ;
        RECT 0.000 2049.515 2889.180 2052.245 ;
        RECT 0.000 2049.465 462.565 2049.515 ;
        RECT 0.000 2046.805 18.665 2046.855 ;
        RECT 0.000 2044.075 2889.180 2046.805 ;
        RECT 0.000 2044.025 6.705 2044.075 ;
        RECT 0.000 2041.365 91.345 2041.415 ;
        RECT 0.000 2038.635 2889.180 2041.365 ;
        RECT 0.000 2038.585 153.905 2038.635 ;
        RECT 0.000 2035.925 138.725 2035.975 ;
        RECT 0.000 2033.195 2889.180 2035.925 ;
        RECT 0.000 2033.145 206.805 2033.195 ;
        RECT 0.000 2030.485 121.245 2030.535 ;
        RECT 0.000 2027.755 2889.180 2030.485 ;
        RECT 0.000 2027.705 4.865 2027.755 ;
        RECT 0.000 2025.045 107.905 2025.095 ;
        RECT 0.000 2022.315 2889.180 2025.045 ;
        RECT 0.000 2022.265 95.485 2022.315 ;
        RECT 0.000 2019.605 254.185 2019.655 ;
        RECT 0.000 2016.875 2889.180 2019.605 ;
        RECT 0.000 2016.825 13.605 2016.875 ;
        RECT 0.000 2014.165 137.805 2014.215 ;
        RECT 0.000 2011.435 2889.180 2014.165 ;
        RECT 0.000 2011.385 32.465 2011.435 ;
        RECT 0.000 2008.725 157.585 2008.775 ;
        RECT 0.000 2005.995 2889.180 2008.725 ;
        RECT 0.000 2005.945 3.945 2005.995 ;
        RECT 0.000 2003.285 109.285 2003.335 ;
        RECT 0.000 2000.555 2889.180 2003.285 ;
        RECT 0.000 2000.505 29.705 2000.555 ;
        RECT 0.000 1997.845 36.145 1997.895 ;
        RECT 0.000 1995.115 2889.180 1997.845 ;
        RECT 0.000 1995.065 50.865 1995.115 ;
        RECT 0.000 1992.405 93.185 1992.455 ;
        RECT 0.000 1989.675 2889.180 1992.405 ;
        RECT 0.000 1989.625 12.685 1989.675 ;
        RECT 0.000 1986.965 48.105 1987.015 ;
        RECT 0.000 1984.235 2889.180 1986.965 ;
        RECT 0.000 1984.185 9.925 1984.235 ;
        RECT 0.000 1981.525 15.905 1981.575 ;
        RECT 0.000 1978.795 2889.180 1981.525 ;
        RECT 0.000 1978.745 32.465 1978.795 ;
        RECT 0.000 1976.085 149.305 1976.135 ;
        RECT 0.000 1973.355 2889.180 1976.085 ;
        RECT 0.000 1973.305 836.545 1973.355 ;
        RECT 0.000 1970.645 65.125 1970.695 ;
        RECT 0.000 1967.915 2889.180 1970.645 ;
        RECT 0.000 1967.865 6.245 1967.915 ;
        RECT 0.000 1965.205 89.505 1965.255 ;
        RECT 0.000 1962.475 2889.180 1965.205 ;
        RECT 0.000 1962.425 21.885 1962.475 ;
        RECT 0.000 1959.765 187.025 1959.815 ;
        RECT 0.000 1957.035 2889.180 1959.765 ;
        RECT 0.000 1956.985 37.525 1957.035 ;
        RECT 0.000 1954.325 173.225 1954.375 ;
        RECT 0.000 1951.595 2889.180 1954.325 ;
        RECT 0.000 1951.545 50.865 1951.595 ;
        RECT 0.000 1948.885 6.705 1948.935 ;
        RECT 0.000 1946.155 2889.180 1948.885 ;
        RECT 0.000 1946.105 71.105 1946.155 ;
        RECT 0.000 1943.445 22.345 1943.495 ;
        RECT 0.000 1940.715 2889.180 1943.445 ;
        RECT 0.000 1940.665 39.825 1940.715 ;
        RECT 0.000 1938.005 186.105 1938.055 ;
        RECT 0.000 1935.275 2889.180 1938.005 ;
        RECT 0.000 1935.225 93.645 1935.275 ;
        RECT 0.000 1932.565 373.785 1932.615 ;
        RECT 0.000 1929.835 2889.180 1932.565 ;
        RECT 0.000 1929.785 65.125 1929.835 ;
        RECT 0.000 1927.125 6.245 1927.175 ;
        RECT 0.000 1924.395 2889.180 1927.125 ;
        RECT 0.000 1924.345 191.165 1924.395 ;
        RECT 0.000 1921.685 140.105 1921.735 ;
        RECT 0.000 1918.955 2889.180 1921.685 ;
        RECT 0.000 1918.905 12.685 1918.955 ;
        RECT 0.000 1916.245 93.185 1916.295 ;
        RECT 0.000 1913.515 2889.180 1916.245 ;
        RECT 0.000 1913.465 318.585 1913.515 ;
        RECT 0.000 1910.805 65.125 1910.855 ;
        RECT 0.000 1908.075 2889.180 1910.805 ;
        RECT 0.000 1908.025 50.405 1908.075 ;
        RECT 0.000 1905.365 371.945 1905.415 ;
        RECT 0.000 1902.635 2889.180 1905.365 ;
        RECT 0.000 1902.585 245.445 1902.635 ;
        RECT 0.000 1899.925 43.965 1899.975 ;
        RECT 0.000 1897.195 2889.180 1899.925 ;
        RECT 0.000 1897.145 122.165 1897.195 ;
        RECT 0.000 1894.485 64.665 1894.535 ;
        RECT 0.000 1891.755 2889.180 1894.485 ;
        RECT 0.000 1891.705 10.845 1891.755 ;
        RECT 0.000 1889.045 105.145 1889.095 ;
        RECT 0.000 1886.315 2889.180 1889.045 ;
        RECT 0.000 1886.265 207.725 1886.315 ;
        RECT 0.000 1883.605 46.725 1883.655 ;
        RECT 0.000 1880.875 2889.180 1883.605 ;
        RECT 0.000 1880.825 17.745 1880.875 ;
        RECT 0.000 1878.165 24.645 1878.215 ;
        RECT 0.000 1875.435 2889.180 1878.165 ;
        RECT 0.000 1875.385 153.445 1875.435 ;
        RECT 0.000 1872.725 241.305 1872.775 ;
        RECT 0.000 1869.995 2889.180 1872.725 ;
        RECT 0.000 1869.945 94.565 1869.995 ;
        RECT 0.000 1867.285 30.165 1867.335 ;
        RECT 0.000 1864.555 2889.180 1867.285 ;
        RECT 0.000 1864.505 37.065 1864.555 ;
        RECT 0.000 1861.845 53.625 1861.895 ;
        RECT 0.000 1859.115 2889.180 1861.845 ;
        RECT 0.000 1859.065 348.025 1859.115 ;
        RECT 0.000 1856.405 164.025 1856.455 ;
        RECT 0.000 1853.675 2889.180 1856.405 ;
        RECT 0.000 1853.625 178.745 1853.675 ;
        RECT 0.000 1850.965 93.185 1851.015 ;
        RECT 0.000 1848.235 2889.180 1850.965 ;
        RECT 0.000 1848.185 15.445 1848.235 ;
        RECT 0.000 1845.525 15.905 1845.575 ;
        RECT 0.000 1842.795 2889.180 1845.525 ;
        RECT 0.000 1842.745 39.825 1842.795 ;
        RECT 0.000 1840.085 77.545 1840.135 ;
        RECT 0.000 1837.355 2889.180 1840.085 ;
        RECT 0.000 1837.305 22.805 1837.355 ;
        RECT 0.000 1834.645 19.585 1834.695 ;
        RECT 0.000 1831.915 2889.180 1834.645 ;
        RECT 0.000 1831.865 177.365 1831.915 ;
        RECT 0.000 1829.205 37.065 1829.255 ;
        RECT 0.000 1826.475 2889.180 1829.205 ;
        RECT 0.000 1826.425 160.805 1826.475 ;
        RECT 0.000 1823.765 15.905 1823.815 ;
        RECT 0.000 1821.035 2889.180 1823.765 ;
        RECT 0.000 1820.985 85.825 1821.035 ;
        RECT 0.000 1818.325 133.665 1818.375 ;
        RECT 0.000 1815.595 2889.180 1818.325 ;
        RECT 0.000 1815.545 554.565 1815.595 ;
        RECT 0.000 1812.885 22.345 1812.935 ;
        RECT 0.000 1810.155 2889.180 1812.885 ;
        RECT 0.000 1810.105 15.445 1810.155 ;
        RECT 0.000 1807.445 81.685 1807.495 ;
        RECT 0.000 1804.715 2889.180 1807.445 ;
        RECT 0.000 1804.665 163.105 1804.715 ;
        RECT 0.000 1802.005 141.025 1802.055 ;
        RECT 0.000 1799.275 2889.180 1802.005 ;
        RECT 0.000 1799.225 384.365 1799.275 ;
        RECT 0.000 1796.565 7.625 1796.615 ;
        RECT 0.000 1793.835 2889.180 1796.565 ;
        RECT 0.000 1793.785 328.245 1793.835 ;
        RECT 0.000 1791.125 23.265 1791.175 ;
        RECT 0.000 1788.395 2889.180 1791.125 ;
        RECT 0.000 1788.345 50.865 1788.395 ;
        RECT 0.000 1785.685 37.065 1785.735 ;
        RECT 0.000 1782.955 2889.180 1785.685 ;
        RECT 0.000 1782.905 170.465 1782.955 ;
        RECT 0.000 1780.245 111.125 1780.295 ;
        RECT 0.000 1777.515 2889.180 1780.245 ;
        RECT 0.000 1777.465 384.825 1777.515 ;
        RECT 0.000 1774.805 429.905 1774.855 ;
        RECT 0.000 1772.075 2889.180 1774.805 ;
        RECT 0.000 1772.025 331.465 1772.075 ;
        RECT 0.000 1769.365 528.805 1769.415 ;
        RECT 0.000 1766.635 2889.180 1769.365 ;
        RECT 0.000 1766.585 303.405 1766.635 ;
        RECT 0.000 1763.925 539.385 1763.975 ;
        RECT 0.000 1761.195 2889.180 1763.925 ;
        RECT 0.000 1761.145 317.665 1761.195 ;
        RECT 0.000 1758.485 338.365 1758.535 ;
        RECT 0.000 1755.755 2889.180 1758.485 ;
        RECT 0.000 1755.705 21.425 1755.755 ;
        RECT 0.000 1753.045 1046.305 1753.095 ;
        RECT 0.000 1750.315 2889.180 1753.045 ;
        RECT 0.000 1750.265 115.265 1750.315 ;
        RECT 0.000 1747.605 15.905 1747.655 ;
        RECT 0.000 1744.875 2889.180 1747.605 ;
        RECT 0.000 1744.825 59.145 1744.875 ;
        RECT 0.000 1742.165 43.965 1742.215 ;
        RECT 0.000 1739.435 2889.180 1742.165 ;
        RECT 0.000 1739.385 181.045 1739.435 ;
        RECT 0.000 1736.725 171.845 1736.775 ;
        RECT 0.000 1733.995 2889.180 1736.725 ;
        RECT 0.000 1733.945 217.845 1733.995 ;
        RECT 0.000 1731.285 168.625 1731.335 ;
        RECT 0.000 1728.555 2889.180 1731.285 ;
        RECT 0.000 1728.505 21.425 1728.555 ;
        RECT 0.000 1725.845 15.905 1725.895 ;
        RECT 0.000 1723.115 2889.180 1725.845 ;
        RECT 0.000 1723.065 163.105 1723.115 ;
        RECT 0.000 1720.405 64.665 1720.455 ;
        RECT 0.000 1717.675 2889.180 1720.405 ;
        RECT 0.000 1717.625 190.245 1717.675 ;
        RECT 0.000 1714.965 49.485 1715.015 ;
        RECT 0.000 1712.235 2889.180 1714.965 ;
        RECT 0.000 1712.185 34.305 1712.235 ;
        RECT 0.000 1709.525 62.365 1709.575 ;
        RECT 0.000 1706.795 2889.180 1709.525 ;
        RECT 0.000 1706.745 19.585 1706.795 ;
        RECT 0.000 1704.085 91.805 1704.135 ;
        RECT 0.000 1701.355 2889.180 1704.085 ;
        RECT 0.000 1701.305 149.765 1701.355 ;
        RECT 0.000 1698.645 138.725 1698.695 ;
        RECT 0.000 1695.915 2889.180 1698.645 ;
        RECT 0.000 1695.865 425.765 1695.915 ;
        RECT 0.000 1693.205 16.825 1693.255 ;
        RECT 0.000 1690.475 2889.180 1693.205 ;
        RECT 0.000 1690.425 106.985 1690.475 ;
        RECT 0.000 1687.765 60.065 1687.815 ;
        RECT 0.000 1685.035 2889.180 1687.765 ;
        RECT 0.000 1684.985 78.925 1685.035 ;
        RECT 0.000 1682.325 43.965 1682.375 ;
        RECT 0.000 1679.595 2889.180 1682.325 ;
        RECT 0.000 1679.545 323.185 1679.595 ;
        RECT 0.000 1676.885 57.765 1676.935 ;
        RECT 0.000 1674.155 2889.180 1676.885 ;
        RECT 0.000 1674.105 183.345 1674.155 ;
        RECT 0.000 1671.445 16.825 1671.495 ;
        RECT 0.000 1668.715 2889.180 1671.445 ;
        RECT 0.000 1668.665 144.245 1668.715 ;
        RECT 0.000 1666.005 214.165 1666.055 ;
        RECT 0.000 1663.275 2889.180 1666.005 ;
        RECT 0.000 1663.225 41.665 1663.275 ;
        RECT 0.000 1660.565 72.025 1660.615 ;
        RECT 0.000 1657.835 2889.180 1660.565 ;
        RECT 0.000 1657.785 115.725 1657.835 ;
        RECT 0.000 1655.125 17.285 1655.175 ;
        RECT 0.000 1652.395 2889.180 1655.125 ;
        RECT 0.000 1652.345 212.325 1652.395 ;
        RECT 0.000 1649.685 324.565 1649.735 ;
        RECT 0.000 1646.955 2889.180 1649.685 ;
        RECT 0.000 1646.905 37.985 1646.955 ;
        RECT 0.000 1644.245 225.665 1644.295 ;
        RECT 0.000 1641.515 2889.180 1644.245 ;
        RECT 0.000 1641.465 113.885 1641.515 ;
        RECT 0.000 1638.805 26.945 1638.855 ;
        RECT 0.000 1636.075 2889.180 1638.805 ;
        RECT 0.000 1636.025 16.825 1636.075 ;
        RECT 0.000 1633.365 51.325 1633.415 ;
        RECT 0.000 1630.635 2889.180 1633.365 ;
        RECT 0.000 1630.585 20.965 1630.635 ;
        RECT 0.000 1627.925 31.545 1627.975 ;
        RECT 0.000 1625.195 2889.180 1627.925 ;
        RECT 0.000 1625.145 88.585 1625.195 ;
        RECT 0.000 1622.485 1926.285 1622.535 ;
        RECT 0.000 1619.755 2889.180 1622.485 ;
        RECT 0.000 1619.705 191.165 1619.755 ;
        RECT 0.000 1617.045 129.525 1617.095 ;
        RECT 0.000 1614.315 2889.180 1617.045 ;
        RECT 0.000 1614.265 20.965 1614.315 ;
        RECT 0.000 1611.605 47.645 1611.655 ;
        RECT 0.000 1608.875 2889.180 1611.605 ;
        RECT 0.000 1608.825 239.465 1608.875 ;
        RECT 0.000 1606.165 35.685 1606.215 ;
        RECT 0.000 1603.435 2889.180 1606.165 ;
        RECT 0.000 1603.385 20.965 1603.435 ;
        RECT 0.000 1600.725 92.725 1600.775 ;
        RECT 0.000 1597.995 2889.180 1600.725 ;
        RECT 0.000 1597.945 116.185 1597.995 ;
        RECT 0.000 1595.285 486.025 1595.335 ;
        RECT 0.000 1592.555 2889.180 1595.285 ;
        RECT 0.000 1592.505 141.945 1592.555 ;
        RECT 0.000 1589.845 33.845 1589.895 ;
        RECT 0.000 1587.115 2889.180 1589.845 ;
        RECT 0.000 1587.065 19.125 1587.115 ;
        RECT 0.000 1584.405 172.305 1584.455 ;
        RECT 0.000 1581.675 2889.180 1584.405 ;
        RECT 0.000 1581.625 49.485 1581.675 ;
        RECT 0.000 1578.965 75.705 1579.015 ;
        RECT 0.000 1576.235 2889.180 1578.965 ;
        RECT 0.000 1576.185 155.745 1576.235 ;
        RECT 0.000 1573.525 144.705 1573.575 ;
        RECT 0.000 1570.795 2889.180 1573.525 ;
        RECT 0.000 1570.745 300.185 1570.795 ;
        RECT 0.000 1568.085 23.265 1568.135 ;
        RECT 0.000 1565.355 2889.180 1568.085 ;
        RECT 0.000 1565.305 113.885 1565.355 ;
        RECT 0.000 1562.645 63.285 1562.695 ;
        RECT 0.000 1559.915 2889.180 1562.645 ;
        RECT 0.000 1559.865 149.765 1559.915 ;
        RECT 0.000 1557.205 77.085 1557.255 ;
        RECT 0.000 1554.475 2889.180 1557.205 ;
        RECT 0.000 1554.425 20.965 1554.475 ;
        RECT 0.000 1551.765 60.065 1551.815 ;
        RECT 0.000 1549.035 2889.180 1551.765 ;
        RECT 0.000 1548.985 160.345 1549.035 ;
        RECT 0.000 1546.325 120.785 1546.375 ;
        RECT 0.000 1543.595 2889.180 1546.325 ;
        RECT 0.000 1543.545 359.525 1543.595 ;
        RECT 0.000 1540.885 411.965 1540.935 ;
        RECT 0.000 1538.155 2889.180 1540.885 ;
        RECT 0.000 1538.105 94.565 1538.155 ;
        RECT 0.000 1535.445 32.925 1535.495 ;
        RECT 0.000 1532.715 2889.180 1535.445 ;
        RECT 0.000 1532.665 17.285 1532.715 ;
        RECT 0.000 1530.005 79.385 1530.055 ;
        RECT 0.000 1527.275 2889.180 1530.005 ;
        RECT 0.000 1527.225 155.745 1527.275 ;
        RECT 0.000 1524.565 156.205 1524.615 ;
        RECT 0.000 1521.835 2889.180 1524.565 ;
        RECT 0.000 1521.785 20.505 1521.835 ;
        RECT 0.000 1519.125 33.385 1519.175 ;
        RECT 0.000 1516.395 2889.180 1519.125 ;
        RECT 0.000 1516.345 65.125 1516.395 ;
        RECT 0.000 1513.685 108.365 1513.735 ;
        RECT 0.000 1510.955 2889.180 1513.685 ;
        RECT 0.000 1510.905 422.545 1510.955 ;
        RECT 0.000 1508.245 79.385 1508.295 ;
        RECT 0.000 1505.515 2889.180 1508.245 ;
        RECT 0.000 1505.465 122.625 1505.515 ;
        RECT 0.000 1502.805 51.325 1502.855 ;
        RECT 0.000 1500.075 2889.180 1502.805 ;
        RECT 0.000 1500.025 450.605 1500.075 ;
        RECT 0.000 1497.365 65.125 1497.415 ;
        RECT 0.000 1494.635 2889.180 1497.365 ;
        RECT 0.000 1494.585 32.465 1494.635 ;
        RECT 0.000 1491.925 50.405 1491.975 ;
        RECT 0.000 1489.195 2889.180 1491.925 ;
        RECT 0.000 1489.145 163.105 1489.195 ;
        RECT 0.000 1486.485 26.485 1486.535 ;
        RECT 0.000 1483.755 2889.180 1486.485 ;
        RECT 0.000 1483.705 95.485 1483.755 ;
        RECT 0.000 1481.045 72.025 1481.095 ;
        RECT 0.000 1478.315 2889.180 1481.045 ;
        RECT 0.000 1478.265 170.005 1478.315 ;
        RECT 0.000 1475.605 47.645 1475.655 ;
        RECT 0.000 1472.875 2889.180 1475.605 ;
        RECT 0.000 1472.825 20.045 1472.875 ;
        RECT 0.000 1470.165 111.125 1470.215 ;
        RECT 0.000 1467.435 2889.180 1470.165 ;
        RECT 0.000 1467.385 183.345 1467.435 ;
        RECT 0.000 1464.725 333.765 1464.775 ;
        RECT 0.000 1461.995 2889.180 1464.725 ;
        RECT 0.000 1461.945 89.045 1461.995 ;
        RECT 0.000 1459.285 65.125 1459.335 ;
        RECT 0.000 1456.555 2889.180 1459.285 ;
        RECT 0.000 1456.505 117.105 1456.555 ;
        RECT 0.000 1453.845 57.305 1453.895 ;
        RECT 0.000 1451.115 2889.180 1453.845 ;
        RECT 0.000 1451.065 97.785 1451.115 ;
        RECT 0.000 1448.405 570.205 1448.455 ;
        RECT 0.000 1445.675 2889.180 1448.405 ;
        RECT 0.000 1445.625 325.025 1445.675 ;
        RECT 0.000 1442.965 333.305 1443.015 ;
        RECT 0.000 1440.235 2889.180 1442.965 ;
        RECT 0.000 1440.185 379.305 1440.235 ;
        RECT 0.000 1437.525 366.425 1437.575 ;
        RECT 0.000 1434.795 2889.180 1437.525 ;
        RECT 0.000 1434.745 353.085 1434.795 ;
        RECT 0.000 1432.085 241.305 1432.135 ;
        RECT 0.000 1429.355 2889.180 1432.085 ;
        RECT 0.000 1429.305 125.385 1429.355 ;
        RECT 0.000 1426.645 46.725 1426.695 ;
        RECT 0.000 1423.915 2889.180 1426.645 ;
        RECT 0.000 1423.865 78.925 1423.915 ;
        RECT 0.000 1421.205 108.825 1421.255 ;
        RECT 0.000 1418.475 2889.180 1421.205 ;
        RECT 0.000 1418.425 143.785 1418.475 ;
        RECT 0.000 1415.765 198.065 1415.815 ;
        RECT 0.000 1413.035 2889.180 1415.765 ;
        RECT 0.000 1412.985 62.365 1413.035 ;
        RECT 0.000 1410.325 494.305 1410.375 ;
        RECT 0.000 1407.595 2889.180 1410.325 ;
        RECT 0.000 1407.545 208.185 1407.595 ;
        RECT 0.000 1404.885 62.825 1404.935 ;
        RECT 0.000 1402.155 2889.180 1404.885 ;
        RECT 0.000 1402.105 30.625 1402.155 ;
        RECT 0.000 1399.445 30.165 1399.495 ;
        RECT 0.000 1396.715 2889.180 1399.445 ;
        RECT 0.000 1396.665 49.945 1396.715 ;
        RECT 0.000 1394.005 247.745 1394.055 ;
        RECT 0.000 1391.275 2889.180 1394.005 ;
        RECT 0.000 1391.225 75.245 1391.275 ;
        RECT 0.000 1388.565 148.845 1388.615 ;
        RECT 0.000 1385.835 2889.180 1388.565 ;
        RECT 0.000 1385.785 58.225 1385.835 ;
        RECT 0.000 1383.125 19.585 1383.175 ;
        RECT 0.000 1380.395 2889.180 1383.125 ;
        RECT 0.000 1380.345 88.585 1380.395 ;
        RECT 0.000 1377.685 121.245 1377.735 ;
        RECT 0.000 1374.955 2889.180 1377.685 ;
        RECT 0.000 1374.905 20.045 1374.955 ;
        RECT 0.000 1372.245 93.185 1372.295 ;
        RECT 0.000 1369.515 2889.180 1372.245 ;
        RECT 0.000 1369.465 43.045 1369.515 ;
        RECT 0.000 1366.805 167.705 1366.855 ;
        RECT 0.000 1364.075 2889.180 1366.805 ;
        RECT 0.000 1364.025 12.225 1364.075 ;
        RECT 0.000 1361.365 57.765 1361.415 ;
        RECT 0.000 1358.635 2889.180 1361.365 ;
        RECT 0.000 1358.585 74.785 1358.635 ;
        RECT 0.000 1355.925 60.065 1355.975 ;
        RECT 0.000 1353.195 2889.180 1355.925 ;
        RECT 0.000 1353.145 211.405 1353.195 ;
        RECT 0.000 1350.485 195.305 1350.535 ;
        RECT 0.000 1347.755 2889.180 1350.485 ;
        RECT 0.000 1347.705 14.065 1347.755 ;
        RECT 0.000 1345.045 149.305 1345.095 ;
        RECT 0.000 1342.315 2889.180 1345.045 ;
        RECT 0.000 1342.265 45.345 1342.315 ;
        RECT 0.000 1339.605 93.185 1339.655 ;
        RECT 0.000 1336.875 2889.180 1339.605 ;
        RECT 0.000 1336.825 289.145 1336.875 ;
        RECT 0.000 1334.165 696.705 1334.215 ;
        RECT 0.000 1331.435 2889.180 1334.165 ;
        RECT 0.000 1331.385 14.525 1331.435 ;
        RECT 0.000 1328.725 352.625 1328.775 ;
        RECT 0.000 1325.995 2889.180 1328.725 ;
        RECT 0.000 1325.945 106.985 1325.995 ;
        RECT 0.000 1323.285 48.565 1323.335 ;
        RECT 0.000 1320.555 2889.180 1323.285 ;
        RECT 0.000 1320.505 273.505 1320.555 ;
        RECT 0.000 1317.845 88.585 1317.895 ;
        RECT 0.000 1315.115 2889.180 1317.845 ;
        RECT 0.000 1315.065 29.705 1315.115 ;
        RECT 0.000 1312.405 345.725 1312.455 ;
        RECT 0.000 1309.675 2889.180 1312.405 ;
        RECT 0.000 1309.625 29.705 1309.675 ;
        RECT 0.000 1306.965 623.105 1307.015 ;
        RECT 0.000 1304.235 2889.180 1306.965 ;
        RECT 0.000 1304.185 518.225 1304.235 ;
        RECT 0.000 1301.525 92.725 1301.575 ;
        RECT 0.000 1298.795 2889.180 1301.525 ;
        RECT 0.000 1298.745 78.925 1298.795 ;
        RECT 0.000 1296.085 130.445 1296.135 ;
        RECT 0.000 1293.355 2889.180 1296.085 ;
        RECT 0.000 1293.305 29.705 1293.355 ;
        RECT 0.000 1290.645 60.525 1290.695 ;
        RECT 0.000 1287.915 2889.180 1290.645 ;
        RECT 0.000 1287.865 19.585 1287.915 ;
        RECT 0.000 1285.205 62.365 1285.255 ;
        RECT 0.000 1282.475 2889.180 1285.205 ;
        RECT 0.000 1282.425 200.365 1282.475 ;
        RECT 0.000 1279.765 146.545 1279.815 ;
        RECT 0.000 1277.035 2889.180 1279.765 ;
        RECT 0.000 1276.985 44.885 1277.035 ;
        RECT 0.000 1274.325 72.025 1274.375 ;
        RECT 0.000 1271.595 2889.180 1274.325 ;
        RECT 0.000 1271.545 78.465 1271.595 ;
        RECT 0.000 1268.885 26.485 1268.935 ;
        RECT 0.000 1266.155 2889.180 1268.885 ;
        RECT 0.000 1266.105 40.745 1266.155 ;
        RECT 0.000 1263.445 212.325 1263.495 ;
        RECT 0.000 1260.715 2889.180 1263.445 ;
        RECT 0.000 1260.665 66.965 1260.715 ;
        RECT 0.000 1258.005 118.485 1258.055 ;
        RECT 0.000 1255.275 2889.180 1258.005 ;
        RECT 0.000 1255.225 85.825 1255.275 ;
        RECT 0.000 1252.565 247.745 1252.615 ;
        RECT 0.000 1249.835 2889.180 1252.565 ;
        RECT 0.000 1249.785 12.685 1249.835 ;
        RECT 0.000 1247.125 27.865 1247.175 ;
        RECT 0.000 1244.395 2889.180 1247.125 ;
        RECT 0.000 1244.345 201.745 1244.395 ;
        RECT 0.000 1241.685 296.505 1241.735 ;
        RECT 0.000 1238.955 2889.180 1241.685 ;
        RECT 0.000 1238.905 78.925 1238.955 ;
        RECT 0.000 1236.245 219.685 1236.295 ;
        RECT 0.000 1233.515 2889.180 1236.245 ;
        RECT 0.000 1233.465 94.565 1233.515 ;
        RECT 0.000 1230.805 52.705 1230.855 ;
        RECT 0.000 1228.075 2889.180 1230.805 ;
        RECT 0.000 1228.025 75.245 1228.075 ;
        RECT 0.000 1225.365 19.125 1225.415 ;
        RECT 0.000 1222.635 2889.180 1225.365 ;
        RECT 0.000 1222.585 161.725 1222.635 ;
        RECT 0.000 1219.925 80.305 1219.975 ;
        RECT 0.000 1217.195 2889.180 1219.925 ;
        RECT 0.000 1217.145 22.805 1217.195 ;
        RECT 0.000 1214.485 240.845 1214.535 ;
        RECT 0.000 1211.755 2889.180 1214.485 ;
        RECT 0.000 1211.705 135.045 1211.755 ;
        RECT 0.000 1209.045 52.705 1209.095 ;
        RECT 0.000 1206.315 2889.180 1209.045 ;
        RECT 0.000 1206.265 74.325 1206.315 ;
        RECT 0.000 1203.605 33.845 1203.655 ;
        RECT 0.000 1200.875 2889.180 1203.605 ;
        RECT 0.000 1200.825 93.645 1200.875 ;
        RECT 0.000 1198.165 121.245 1198.215 ;
        RECT 0.000 1195.435 2889.180 1198.165 ;
        RECT 0.000 1195.385 15.905 1195.435 ;
        RECT 0.000 1192.725 138.265 1192.775 ;
        RECT 0.000 1189.995 2889.180 1192.725 ;
        RECT 0.000 1189.945 66.505 1189.995 ;
        RECT 0.000 1187.285 46.725 1187.335 ;
        RECT 0.000 1184.555 2889.180 1187.285 ;
        RECT 0.000 1184.505 14.525 1184.555 ;
        RECT 0.000 1181.845 141.945 1181.895 ;
        RECT 0.000 1179.115 2889.180 1181.845 ;
        RECT 0.000 1179.065 347.565 1179.115 ;
        RECT 0.000 1176.405 198.985 1176.455 ;
        RECT 0.000 1173.675 2889.180 1176.405 ;
        RECT 0.000 1173.625 198.065 1173.675 ;
        RECT 0.000 1170.965 72.025 1171.015 ;
        RECT 0.000 1168.235 2889.180 1170.965 ;
        RECT 0.000 1168.185 259.705 1168.235 ;
        RECT 0.000 1165.525 243.145 1165.575 ;
        RECT 0.000 1162.795 2889.180 1165.525 ;
        RECT 0.000 1162.745 22.345 1162.795 ;
        RECT 0.000 1160.085 55.925 1160.135 ;
        RECT 0.000 1157.355 2889.180 1160.085 ;
        RECT 0.000 1157.305 258.325 1157.355 ;
        RECT 0.000 1154.645 110.665 1154.695 ;
        RECT 0.000 1151.915 2889.180 1154.645 ;
        RECT 0.000 1151.865 480.045 1151.915 ;
        RECT 0.000 1149.205 429.905 1149.255 ;
        RECT 0.000 1146.475 2889.180 1149.205 ;
        RECT 0.000 1146.425 424.845 1146.475 ;
        RECT 0.000 1143.765 380.685 1143.815 ;
        RECT 0.000 1141.035 2889.180 1143.765 ;
        RECT 0.000 1140.985 339.285 1141.035 ;
        RECT 0.000 1138.325 82.605 1138.375 ;
        RECT 0.000 1135.595 2889.180 1138.325 ;
        RECT 0.000 1135.545 175.525 1135.595 ;
        RECT 0.000 1132.885 113.425 1132.935 ;
        RECT 0.000 1130.155 2889.180 1132.885 ;
        RECT 0.000 1130.105 37.985 1130.155 ;
        RECT 0.000 1127.445 8.085 1127.495 ;
        RECT 0.000 1124.715 2889.180 1127.445 ;
        RECT 0.000 1124.665 22.345 1124.715 ;
        RECT 0.000 1122.005 689.345 1122.055 ;
        RECT 0.000 1119.275 2889.180 1122.005 ;
        RECT 0.000 1119.225 50.865 1119.275 ;
        RECT 0.000 1116.565 149.305 1116.615 ;
        RECT 0.000 1113.835 2889.180 1116.565 ;
        RECT 0.000 1113.785 22.345 1113.835 ;
        RECT 0.000 1111.125 100.085 1111.175 ;
        RECT 0.000 1108.395 2889.180 1111.125 ;
        RECT 0.000 1108.345 178.745 1108.395 ;
        RECT 0.000 1105.685 52.705 1105.735 ;
        RECT 0.000 1102.955 2889.180 1105.685 ;
        RECT 0.000 1102.905 10.385 1102.955 ;
        RECT 0.000 1100.245 20.965 1100.295 ;
        RECT 0.000 1097.515 2889.180 1100.245 ;
        RECT 0.000 1097.465 134.125 1097.515 ;
        RECT 0.000 1094.805 9.005 1094.855 ;
        RECT 0.000 1092.075 2889.180 1094.805 ;
        RECT 0.000 1092.025 355.385 1092.075 ;
        RECT 0.000 1089.365 77.085 1089.415 ;
        RECT 0.000 1086.635 2889.180 1089.365 ;
        RECT 0.000 1086.585 46.725 1086.635 ;
        RECT 0.000 1083.925 149.305 1083.975 ;
        RECT 0.000 1081.195 2889.180 1083.925 ;
        RECT 0.000 1081.145 215.085 1081.195 ;
        RECT 0.000 1078.485 9.005 1078.535 ;
        RECT 0.000 1075.755 2889.180 1078.485 ;
        RECT 0.000 1075.705 205.425 1075.755 ;
        RECT 0.000 1073.045 56.385 1073.095 ;
        RECT 0.000 1070.315 2889.180 1073.045 ;
        RECT 0.000 1070.265 78.005 1070.315 ;
        RECT 0.000 1067.605 29.705 1067.655 ;
        RECT 0.000 1064.875 2889.180 1067.605 ;
        RECT 0.000 1064.825 387.585 1064.875 ;
        RECT 0.000 1062.165 43.965 1062.215 ;
        RECT 0.000 1059.435 2889.180 1062.165 ;
        RECT 0.000 1059.385 141.945 1059.435 ;
        RECT 0.000 1056.725 82.145 1056.775 ;
        RECT 0.000 1053.995 2889.180 1056.725 ;
        RECT 0.000 1053.945 50.865 1053.995 ;
        RECT 0.000 1051.285 37.065 1051.335 ;
        RECT 0.000 1048.555 2889.180 1051.285 ;
        RECT 0.000 1048.505 6.245 1048.555 ;
        RECT 0.000 1045.845 147.005 1045.895 ;
        RECT 0.000 1043.115 2889.180 1045.845 ;
        RECT 0.000 1043.065 77.085 1043.115 ;
        RECT 0.000 1040.405 26.945 1040.455 ;
        RECT 0.000 1037.675 2889.180 1040.405 ;
        RECT 0.000 1037.625 65.585 1037.675 ;
        RECT 0.000 1034.965 7.165 1035.015 ;
        RECT 0.000 1032.235 2889.180 1034.965 ;
        RECT 0.000 1032.185 113.885 1032.235 ;
        RECT 0.000 1029.525 77.085 1029.575 ;
        RECT 0.000 1026.795 2889.180 1029.525 ;
        RECT 0.000 1026.745 543.065 1026.795 ;
        RECT 0.000 1024.085 145.625 1024.135 ;
        RECT 0.000 1021.355 2889.180 1024.085 ;
        RECT 0.000 1021.305 69.265 1021.355 ;
        RECT 0.000 1018.645 8.085 1018.695 ;
        RECT 0.000 1015.915 2889.180 1018.645 ;
        RECT 0.000 1015.865 46.725 1015.915 ;
        RECT 0.000 1013.205 23.725 1013.255 ;
        RECT 0.000 1010.475 2889.180 1013.205 ;
        RECT 0.000 1010.425 183.345 1010.475 ;
        RECT 0.000 1007.765 9.005 1007.815 ;
        RECT 0.000 1005.035 2889.180 1007.765 ;
        RECT 0.000 1004.985 152.985 1005.035 ;
        RECT 0.000 1002.325 204.505 1002.375 ;
        RECT 0.000 999.595 2889.180 1002.325 ;
        RECT 0.000 999.545 70.645 999.595 ;
        RECT 0.000 996.885 55.465 996.935 ;
        RECT 0.000 994.155 2889.180 996.885 ;
        RECT 0.000 994.105 39.365 994.155 ;
        RECT 0.000 991.445 23.725 991.495 ;
        RECT 0.000 988.715 2889.180 991.445 ;
        RECT 0.000 988.665 234.865 988.715 ;
        RECT 0.000 986.005 197.145 986.055 ;
        RECT 0.000 983.275 2889.180 986.005 ;
        RECT 0.000 983.225 415.185 983.275 ;
        RECT 0.000 980.565 7.625 980.615 ;
        RECT 0.000 977.835 2889.180 980.565 ;
        RECT 0.000 977.785 69.725 977.835 ;
        RECT 0.000 975.125 212.325 975.175 ;
        RECT 0.000 972.395 2889.180 975.125 ;
        RECT 0.000 972.345 40.745 972.395 ;
        RECT 0.000 969.685 8.545 969.735 ;
        RECT 0.000 966.955 2889.180 969.685 ;
        RECT 0.000 966.905 85.825 966.955 ;
        RECT 0.000 964.245 184.265 964.295 ;
        RECT 0.000 961.515 2889.180 964.245 ;
        RECT 0.000 961.465 6.705 961.515 ;
        RECT 0.000 958.805 85.825 958.855 ;
        RECT 0.000 956.075 2889.180 958.805 ;
        RECT 0.000 956.025 219.225 956.075 ;
        RECT 0.000 953.365 58.225 953.415 ;
        RECT 0.000 950.635 2889.180 953.365 ;
        RECT 0.000 950.585 22.805 950.635 ;
        RECT 0.000 947.925 241.765 947.975 ;
        RECT 0.000 945.195 2889.180 947.925 ;
        RECT 0.000 945.145 515.465 945.195 ;
        RECT 0.000 942.485 17.285 942.535 ;
        RECT 0.000 939.755 2889.180 942.485 ;
        RECT 0.000 939.705 86.745 939.755 ;
        RECT 0.000 937.045 55.465 937.095 ;
        RECT 0.000 934.315 2889.180 937.045 ;
        RECT 0.000 934.265 370.105 934.315 ;
        RECT 0.000 931.605 9.005 931.655 ;
        RECT 0.000 928.875 2889.180 931.605 ;
        RECT 0.000 928.825 38.905 928.875 ;
        RECT 0.000 926.165 168.165 926.215 ;
        RECT 0.000 923.435 2889.180 926.165 ;
        RECT 0.000 923.385 387.125 923.435 ;
        RECT 0.000 920.725 52.245 920.775 ;
        RECT 0.000 917.995 2889.180 920.725 ;
        RECT 0.000 917.945 78.925 917.995 ;
        RECT 0.000 915.285 16.365 915.335 ;
        RECT 0.000 912.555 2889.180 915.285 ;
        RECT 0.000 912.505 123.085 912.555 ;
        RECT 0.000 909.845 373.325 909.895 ;
        RECT 0.000 907.115 2889.180 909.845 ;
        RECT 0.000 907.065 50.865 907.115 ;
        RECT 0.000 904.405 104.685 904.455 ;
        RECT 0.000 901.675 2889.180 904.405 ;
        RECT 0.000 901.625 8.085 901.675 ;
        RECT 0.000 898.965 34.305 899.015 ;
        RECT 0.000 896.235 2889.180 898.965 ;
        RECT 0.000 896.185 233.485 896.235 ;
        RECT 0.000 893.525 81.685 893.575 ;
        RECT 0.000 890.795 2889.180 893.525 ;
        RECT 0.000 890.745 191.165 890.795 ;
        RECT 0.000 888.085 65.125 888.135 ;
        RECT 0.000 885.355 2889.180 888.085 ;
        RECT 0.000 885.305 48.565 885.355 ;
        RECT 0.000 882.645 18.205 882.695 ;
        RECT 0.000 879.915 2889.180 882.645 ;
        RECT 0.000 879.865 85.825 879.915 ;
        RECT 0.000 877.205 101.005 877.255 ;
        RECT 0.000 874.475 2889.180 877.205 ;
        RECT 0.000 874.425 148.385 874.475 ;
        RECT 0.000 871.765 203.585 871.815 ;
        RECT 0.000 869.035 2889.180 871.765 ;
        RECT 0.000 868.985 441.865 869.035 ;
        RECT 0.000 866.325 65.125 866.375 ;
        RECT 0.000 863.595 2889.180 866.325 ;
        RECT 0.000 863.545 324.105 863.595 ;
        RECT 0.000 860.885 156.205 860.935 ;
        RECT 0.000 858.155 2889.180 860.885 ;
        RECT 0.000 858.105 114.345 858.155 ;
        RECT 0.000 855.445 83.985 855.495 ;
        RECT 0.000 852.715 2889.180 855.445 ;
        RECT 0.000 852.665 215.545 852.715 ;
        RECT 0.000 850.005 214.165 850.055 ;
        RECT 0.000 847.275 2889.180 850.005 ;
        RECT 0.000 847.225 443.705 847.275 ;
        RECT 0.000 844.565 197.145 844.615 ;
        RECT 0.000 841.835 2889.180 844.565 ;
        RECT 0.000 841.785 254.185 841.835 ;
        RECT 0.000 839.125 303.865 839.175 ;
        RECT 0.000 836.395 2889.180 839.125 ;
        RECT 0.000 836.345 134.125 836.395 ;
        RECT 0.000 833.685 72.485 833.735 ;
        RECT 0.000 830.955 2889.180 833.685 ;
        RECT 0.000 830.905 14.065 830.955 ;
        RECT 0.000 828.245 2.565 828.295 ;
        RECT 0.000 825.515 2889.180 828.245 ;
        RECT 0.000 825.465 29.705 825.515 ;
        RECT 0.000 822.805 139.645 822.855 ;
        RECT 0.000 820.075 2889.180 822.805 ;
        RECT 0.000 820.025 60.065 820.075 ;
        RECT 0.000 817.365 35.225 817.415 ;
        RECT 0.000 814.635 2889.180 817.365 ;
        RECT 0.000 814.585 183.805 814.635 ;
        RECT 0.000 811.925 316.285 811.975 ;
        RECT 0.000 809.195 2889.180 811.925 ;
        RECT 0.000 809.145 49.485 809.195 ;
        RECT 0.000 806.485 213.245 806.535 ;
        RECT 0.000 803.755 2889.180 806.485 ;
        RECT 0.000 803.705 77.545 803.755 ;
        RECT 0.000 801.045 8.545 801.095 ;
        RECT 0.000 798.315 2889.180 801.045 ;
        RECT 0.000 798.265 22.345 798.315 ;
        RECT 0.000 795.605 634.145 795.655 ;
        RECT 0.000 792.875 2889.180 795.605 ;
        RECT 0.000 792.825 178.745 792.875 ;
        RECT 0.000 790.165 164.945 790.215 ;
        RECT 0.000 787.435 2889.180 790.165 ;
        RECT 0.000 787.385 61.445 787.435 ;
        RECT 0.000 784.725 89.505 784.775 ;
        RECT 0.000 781.995 2889.180 784.725 ;
        RECT 0.000 781.945 114.805 781.995 ;
        RECT 0.000 779.285 43.965 779.335 ;
        RECT 0.000 776.555 2889.180 779.285 ;
        RECT 0.000 776.505 42.585 776.555 ;
        RECT 0.000 773.845 9.005 773.895 ;
        RECT 0.000 771.115 2889.180 773.845 ;
        RECT 0.000 771.065 59.145 771.115 ;
        RECT 0.000 768.405 184.725 768.455 ;
        RECT 0.000 765.675 2889.180 768.405 ;
        RECT 0.000 765.625 78.925 765.675 ;
        RECT 0.000 762.965 258.325 763.015 ;
        RECT 0.000 760.235 2889.180 762.965 ;
        RECT 0.000 760.185 15.445 760.235 ;
        RECT 0.000 757.525 3.025 757.575 ;
        RECT 0.000 754.795 2889.180 757.525 ;
        RECT 0.000 754.745 32.925 754.795 ;
        RECT 0.000 752.085 110.665 752.135 ;
        RECT 0.000 749.355 2889.180 752.085 ;
        RECT 0.000 749.305 272.585 749.355 ;
        RECT 0.000 746.645 15.905 746.695 ;
        RECT 0.000 743.915 2889.180 746.645 ;
        RECT 0.000 743.865 94.565 743.915 ;
        RECT 0.000 741.205 65.125 741.255 ;
        RECT 0.000 738.475 2889.180 741.205 ;
        RECT 0.000 738.425 338.365 738.475 ;
        RECT 0.000 735.765 213.245 735.815 ;
        RECT 0.000 733.035 2889.180 735.765 ;
        RECT 0.000 732.985 199.905 733.035 ;
        RECT 0.000 730.325 31.085 730.375 ;
        RECT 0.000 727.595 2889.180 730.325 ;
        RECT 0.000 727.545 761.105 727.595 ;
        RECT 0.000 724.885 148.845 724.935 ;
        RECT 0.000 722.155 2889.180 724.885 ;
        RECT 0.000 722.105 213.705 722.155 ;
        RECT 0.000 719.445 7.625 719.495 ;
        RECT 0.000 716.715 2889.180 719.445 ;
        RECT 0.000 716.665 57.765 716.715 ;
        RECT 0.000 714.005 189.325 714.055 ;
        RECT 0.000 711.275 2889.180 714.005 ;
        RECT 0.000 711.225 14.065 711.275 ;
        RECT 0.000 708.565 43.965 708.615 ;
        RECT 0.000 705.835 2889.180 708.565 ;
        RECT 0.000 705.785 210.485 705.835 ;
        RECT 0.000 703.125 27.865 703.175 ;
        RECT 0.000 700.395 2889.180 703.125 ;
        RECT 0.000 700.345 282.245 700.395 ;
        RECT 0.000 697.685 329.165 697.735 ;
        RECT 0.000 694.955 2889.180 697.685 ;
        RECT 0.000 694.905 12.225 694.955 ;
        RECT 0.000 692.245 43.965 692.295 ;
        RECT 0.000 689.515 2889.180 692.245 ;
        RECT 0.000 689.465 185.185 689.515 ;
        RECT 0.000 686.805 25.565 686.855 ;
        RECT 0.000 684.075 2889.180 686.805 ;
        RECT 0.000 684.025 2.565 684.075 ;
        RECT 0.000 681.365 85.365 681.415 ;
        RECT 0.000 678.635 2889.180 681.365 ;
        RECT 0.000 678.585 70.185 678.635 ;
        RECT 0.000 675.925 280.865 675.975 ;
        RECT 0.000 673.195 2889.180 675.925 ;
        RECT 0.000 673.145 42.585 673.195 ;
        RECT 0.000 670.485 2.565 670.535 ;
        RECT 0.000 667.755 2889.180 670.485 ;
        RECT 0.000 667.705 209.565 667.755 ;
        RECT 0.000 665.045 128.145 665.095 ;
        RECT 0.000 662.315 2889.180 665.045 ;
        RECT 0.000 662.265 14.985 662.315 ;
        RECT 0.000 659.605 15.905 659.655 ;
        RECT 0.000 656.875 2889.180 659.605 ;
        RECT 0.000 656.825 31.085 656.875 ;
        RECT 0.000 654.165 408.745 654.215 ;
        RECT 0.000 651.435 2889.180 654.165 ;
        RECT 0.000 651.385 76.165 651.435 ;
        RECT 0.000 648.725 165.865 648.775 ;
        RECT 0.000 645.995 2889.180 648.725 ;
        RECT 0.000 645.945 2.565 645.995 ;
        RECT 0.000 643.285 57.765 643.335 ;
        RECT 0.000 640.555 2889.180 643.285 ;
        RECT 0.000 640.505 71.105 640.555 ;
        RECT 0.000 637.845 233.025 637.895 ;
        RECT 0.000 635.115 2889.180 637.845 ;
        RECT 0.000 635.065 163.105 635.115 ;
        RECT 0.000 632.405 100.085 632.455 ;
        RECT 0.000 629.675 2889.180 632.405 ;
        RECT 0.000 629.625 183.345 629.675 ;
        RECT 0.000 626.965 467.625 627.015 ;
        RECT 0.000 624.235 2889.180 626.965 ;
        RECT 0.000 624.185 59.605 624.235 ;
        RECT 0.000 621.525 36.605 621.575 ;
        RECT 0.000 618.795 2889.180 621.525 ;
        RECT 0.000 618.745 2.565 618.795 ;
        RECT 0.000 616.085 205.425 616.135 ;
        RECT 0.000 613.355 2889.180 616.085 ;
        RECT 0.000 613.305 97.325 613.355 ;
        RECT 0.000 610.645 45.805 610.695 ;
        RECT 0.000 607.915 2889.180 610.645 ;
        RECT 0.000 607.865 19.125 607.915 ;
        RECT 0.000 605.205 141.025 605.255 ;
        RECT 0.000 602.475 2889.180 605.205 ;
        RECT 0.000 602.425 75.245 602.475 ;
        RECT 0.000 599.765 92.725 599.815 ;
        RECT 0.000 597.035 2889.180 599.765 ;
        RECT 0.000 596.985 191.165 597.035 ;
        RECT 0.000 594.325 57.765 594.375 ;
        RECT 0.000 591.595 2889.180 594.325 ;
        RECT 0.000 591.545 2.565 591.595 ;
        RECT 0.000 588.885 34.765 588.935 ;
        RECT 0.000 586.155 2889.180 588.885 ;
        RECT 0.000 586.105 14.065 586.155 ;
        RECT 0.000 583.445 268.445 583.495 ;
        RECT 0.000 580.715 2889.180 583.445 ;
        RECT 0.000 580.665 331.465 580.715 ;
        RECT 0.000 578.005 16.825 578.055 ;
        RECT 0.000 575.275 2889.180 578.005 ;
        RECT 0.000 575.225 189.785 575.275 ;
        RECT 0.000 572.565 59.145 572.615 ;
        RECT 0.000 569.835 2889.180 572.565 ;
        RECT 0.000 569.785 17.285 569.835 ;
        RECT 0.000 567.125 2.565 567.175 ;
        RECT 0.000 564.395 2889.180 567.125 ;
        RECT 0.000 564.345 123.085 564.395 ;
        RECT 0.000 561.685 44.425 561.735 ;
        RECT 0.000 558.955 2889.180 561.685 ;
        RECT 0.000 558.905 155.745 558.955 ;
        RECT 0.000 556.245 184.265 556.295 ;
        RECT 0.000 553.515 2889.180 556.245 ;
        RECT 0.000 553.465 157.585 553.515 ;
        RECT 0.000 550.805 76.625 550.855 ;
        RECT 0.000 548.075 2889.180 550.805 ;
        RECT 0.000 548.025 50.865 548.075 ;
        RECT 0.000 545.365 136.885 545.415 ;
        RECT 0.000 542.635 2889.180 545.365 ;
        RECT 0.000 542.585 6.705 542.635 ;
        RECT 0.000 539.925 115.265 539.975 ;
        RECT 0.000 537.195 2889.180 539.925 ;
        RECT 0.000 537.145 10.385 537.195 ;
        RECT 0.000 534.485 249.585 534.535 ;
        RECT 0.000 531.755 2889.180 534.485 ;
        RECT 0.000 531.705 40.745 531.755 ;
        RECT 0.000 529.045 287.765 529.095 ;
        RECT 0.000 526.315 2889.180 529.045 ;
        RECT 0.000 526.265 2.565 526.315 ;
        RECT 0.000 523.605 27.865 523.655 ;
        RECT 0.000 520.875 2889.180 523.605 ;
        RECT 0.000 520.825 396.785 520.875 ;
        RECT 0.000 518.165 60.065 518.215 ;
        RECT 0.000 515.435 2889.180 518.165 ;
        RECT 0.000 515.385 12.225 515.435 ;
        RECT 0.000 512.725 54.085 512.775 ;
        RECT 0.000 509.995 2889.180 512.725 ;
        RECT 0.000 509.945 75.245 509.995 ;
        RECT 0.000 507.285 37.065 507.335 ;
        RECT 0.000 504.555 2889.180 507.285 ;
        RECT 0.000 504.505 283.165 504.555 ;
        RECT 0.000 501.845 188.865 501.895 ;
        RECT 0.000 499.115 2889.180 501.845 ;
        RECT 0.000 499.065 2.565 499.115 ;
        RECT 0.000 496.405 36.145 496.455 ;
        RECT 0.000 493.675 2889.180 496.405 ;
        RECT 0.000 493.625 245.445 493.675 ;
        RECT 0.000 490.965 9.005 491.015 ;
        RECT 0.000 488.235 2889.180 490.965 ;
        RECT 0.000 488.185 49.025 488.235 ;
        RECT 0.000 485.525 7.625 485.575 ;
        RECT 0.000 482.795 2889.180 485.525 ;
        RECT 0.000 482.745 71.565 482.795 ;
        RECT 0.000 480.085 232.565 480.135 ;
        RECT 0.000 477.355 2889.180 480.085 ;
        RECT 0.000 477.305 44.425 477.355 ;
        RECT 0.000 474.645 26.485 474.695 ;
        RECT 0.000 471.915 2889.180 474.645 ;
        RECT 0.000 471.865 58.685 471.915 ;
        RECT 0.000 469.205 141.945 469.255 ;
        RECT 0.000 466.475 2889.180 469.205 ;
        RECT 0.000 466.425 113.885 466.475 ;
        RECT 0.000 463.765 193.005 463.815 ;
        RECT 0.000 461.035 2889.180 463.765 ;
        RECT 0.000 460.985 93.645 461.035 ;
        RECT 0.000 458.325 57.305 458.375 ;
        RECT 0.000 455.595 2889.180 458.325 ;
        RECT 0.000 455.545 185.185 455.595 ;
        RECT 0.000 452.885 35.685 452.935 ;
        RECT 0.000 450.155 2889.180 452.885 ;
        RECT 0.000 450.105 37.065 450.155 ;
        RECT 0.000 447.445 2.565 447.495 ;
        RECT 0.000 444.715 2889.180 447.445 ;
        RECT 0.000 444.665 352.625 444.715 ;
        RECT 0.000 442.005 89.045 442.055 ;
        RECT 0.000 439.275 2889.180 442.005 ;
        RECT 0.000 439.225 15.445 439.275 ;
        RECT 0.000 436.565 193.465 436.615 ;
        RECT 0.000 433.835 2889.180 436.565 ;
        RECT 0.000 433.785 114.345 433.835 ;
        RECT 0.000 431.125 475.445 431.175 ;
        RECT 0.000 428.395 2889.180 431.125 ;
        RECT 0.000 428.345 122.165 428.395 ;
        RECT 0.000 425.685 81.685 425.735 ;
        RECT 0.000 422.955 2889.180 425.685 ;
        RECT 0.000 422.905 49.025 422.955 ;
        RECT 0.000 420.245 121.245 420.295 ;
        RECT 0.000 417.515 2889.180 420.245 ;
        RECT 0.000 417.465 2.565 417.515 ;
        RECT 0.000 414.805 205.425 414.855 ;
        RECT 0.000 412.075 2889.180 414.805 ;
        RECT 0.000 412.025 228.885 412.075 ;
        RECT 0.000 409.365 5.785 409.415 ;
        RECT 0.000 406.635 2889.180 409.365 ;
        RECT 0.000 406.585 170.005 406.635 ;
        RECT 0.000 403.925 452.445 403.975 ;
        RECT 0.000 401.195 2889.180 403.925 ;
        RECT 0.000 401.145 113.885 401.195 ;
        RECT 0.000 398.485 44.425 398.535 ;
        RECT 0.000 395.755 2889.180 398.485 ;
        RECT 0.000 395.705 22.805 395.755 ;
        RECT 0.000 393.045 52.245 393.095 ;
        RECT 0.000 390.315 2889.180 393.045 ;
        RECT 0.000 390.265 10.845 390.315 ;
        RECT 0.000 387.605 53.165 387.655 ;
        RECT 0.000 384.875 2889.180 387.605 ;
        RECT 0.000 384.825 2.565 384.875 ;
        RECT 0.000 382.165 59.145 382.215 ;
        RECT 0.000 379.435 2889.180 382.165 ;
        RECT 0.000 379.385 152.525 379.435 ;
        RECT 0.000 376.725 135.505 376.775 ;
        RECT 0.000 373.995 2889.180 376.725 ;
        RECT 0.000 373.945 480.505 373.995 ;
        RECT 0.000 371.285 9.005 371.335 ;
        RECT 0.000 368.555 2889.180 371.285 ;
        RECT 0.000 368.505 8.085 368.555 ;
        RECT 0.000 365.845 110.205 365.895 ;
        RECT 0.000 363.115 2889.180 365.845 ;
        RECT 0.000 363.065 70.645 363.115 ;
        RECT 0.000 360.405 380.685 360.455 ;
        RECT 0.000 357.675 2889.180 360.405 ;
        RECT 0.000 357.625 310.305 357.675 ;
        RECT 0.000 354.965 355.385 355.015 ;
        RECT 0.000 352.235 2889.180 354.965 ;
        RECT 0.000 352.185 68.805 352.235 ;
        RECT 0.000 349.525 177.365 349.575 ;
        RECT 0.000 346.795 2889.180 349.525 ;
        RECT 0.000 346.745 406.445 346.795 ;
        RECT 0.000 344.085 204.505 344.135 ;
        RECT 0.000 341.355 2889.180 344.085 ;
        RECT 0.000 341.305 115.725 341.355 ;
        RECT 0.000 338.645 104.685 338.695 ;
        RECT 0.000 335.915 2889.180 338.645 ;
        RECT 0.000 335.865 88.125 335.915 ;
        RECT 0.000 333.205 196.225 333.255 ;
        RECT 0.000 330.475 2889.180 333.205 ;
        RECT 0.000 330.425 499.825 330.475 ;
        RECT 0.000 327.765 139.185 327.815 ;
        RECT 0.000 325.035 2889.180 327.765 ;
        RECT 0.000 324.985 43.505 325.035 ;
        RECT 0.000 322.325 43.965 322.375 ;
        RECT 0.000 319.595 2889.180 322.325 ;
        RECT 0.000 319.545 113.885 319.595 ;
        RECT 0.000 316.885 51.325 316.935 ;
        RECT 0.000 314.155 2889.180 316.885 ;
        RECT 0.000 314.105 180.585 314.155 ;
        RECT 0.000 311.445 317.205 311.495 ;
        RECT 0.000 308.715 2889.180 311.445 ;
        RECT 0.000 308.665 172.765 308.715 ;
        RECT 0.000 306.005 135.505 306.055 ;
        RECT 0.000 303.275 2889.180 306.005 ;
        RECT 0.000 303.225 152.985 303.275 ;
        RECT 0.000 300.565 102.385 300.615 ;
        RECT 0.000 297.835 2889.180 300.565 ;
        RECT 0.000 297.785 49.025 297.835 ;
        RECT 0.000 295.125 200.825 295.175 ;
        RECT 0.000 292.395 2889.180 295.125 ;
        RECT 0.000 292.345 63.285 292.395 ;
        RECT 0.000 289.685 33.845 289.735 ;
        RECT 0.000 286.955 2889.180 289.685 ;
        RECT 0.000 286.905 121.245 286.955 ;
        RECT 0.000 284.245 371.945 284.295 ;
        RECT 0.000 281.515 2889.180 284.245 ;
        RECT 0.000 281.465 258.325 281.515 ;
        RECT 0.000 278.805 72.025 278.855 ;
        RECT 0.000 276.075 2889.180 278.805 ;
        RECT 0.000 276.025 41.205 276.075 ;
        RECT 0.000 273.365 156.205 273.415 ;
        RECT 0.000 270.635 2889.180 273.365 ;
        RECT 0.000 270.585 37.525 270.635 ;
        RECT 0.000 267.925 201.745 267.975 ;
        RECT 0.000 265.195 2889.180 267.925 ;
        RECT 0.000 265.145 76.625 265.195 ;
        RECT 0.000 262.485 373.785 262.535 ;
        RECT 0.000 259.755 2889.180 262.485 ;
        RECT 0.000 259.705 267.065 259.755 ;
        RECT 0.000 257.045 100.085 257.095 ;
        RECT 0.000 254.315 2889.180 257.045 ;
        RECT 0.000 254.265 114.805 254.315 ;
        RECT 0.000 251.605 51.325 251.655 ;
        RECT 0.000 248.875 2889.180 251.605 ;
        RECT 0.000 248.825 75.705 248.875 ;
        RECT 0.000 246.165 167.245 246.215 ;
        RECT 0.000 243.435 2889.180 246.165 ;
        RECT 0.000 243.385 130.445 243.435 ;
        RECT 0.000 240.725 37.065 240.775 ;
        RECT 0.000 237.995 2889.180 240.725 ;
        RECT 0.000 237.945 283.165 237.995 ;
        RECT 0.000 235.285 93.185 235.335 ;
        RECT 0.000 232.555 2889.180 235.285 ;
        RECT 0.000 232.505 59.605 232.555 ;
        RECT 0.000 229.845 112.045 229.895 ;
        RECT 0.000 227.115 2889.180 229.845 ;
        RECT 0.000 227.065 60.985 227.115 ;
        RECT 0.000 224.405 46.265 224.455 ;
        RECT 0.000 221.675 2889.180 224.405 ;
        RECT 0.000 221.625 180.125 221.675 ;
        RECT 0.000 218.965 112.965 219.015 ;
        RECT 0.000 216.235 2889.180 218.965 ;
        RECT 0.000 216.185 37.065 216.235 ;
        RECT 0.000 213.525 983.745 213.575 ;
        RECT 0.000 210.795 2889.180 213.525 ;
        RECT 0.000 210.745 65.585 210.795 ;
        RECT 0.000 208.085 101.005 208.135 ;
        RECT 0.000 205.355 2889.180 208.085 ;
        RECT 0.000 205.305 86.745 205.355 ;
        RECT 0.000 202.645 90.425 202.695 ;
        RECT 0.000 199.915 2889.180 202.645 ;
        RECT 0.000 199.865 37.065 199.915 ;
        RECT 0.000 197.205 52.705 197.255 ;
        RECT 0.000 194.475 2889.180 197.205 ;
        RECT 0.000 194.425 104.225 194.475 ;
        RECT 0.000 191.765 52.705 191.815 ;
        RECT 0.000 189.035 2889.180 191.765 ;
        RECT 0.000 188.985 239.465 189.035 ;
        RECT 0.000 186.325 79.385 186.375 ;
        RECT 0.000 183.595 2889.180 186.325 ;
        RECT 0.000 183.545 338.365 183.595 ;
        RECT 0.000 180.885 63.285 180.935 ;
        RECT 0.000 178.155 2889.180 180.885 ;
        RECT 0.000 178.105 317.665 178.155 ;
        RECT 0.000 175.445 113.425 175.495 ;
        RECT 0.000 172.715 2889.180 175.445 ;
        RECT 0.000 172.665 254.185 172.715 ;
        RECT 0.000 170.005 176.445 170.055 ;
        RECT 0.000 167.275 2889.180 170.005 ;
        RECT 0.000 167.225 198.065 167.275 ;
        RECT 0.000 164.565 100.085 164.615 ;
        RECT 0.000 161.835 2889.180 164.565 ;
        RECT 0.000 161.785 159.885 161.835 ;
        RECT 0.000 159.125 88.125 159.175 ;
        RECT 0.000 156.395 2889.180 159.125 ;
        RECT 0.000 156.345 39.825 156.395 ;
        RECT 0.000 153.685 195.305 153.735 ;
        RECT 0.000 150.955 2889.180 153.685 ;
        RECT 0.000 150.905 254.185 150.955 ;
        RECT 0.000 148.245 217.385 148.295 ;
        RECT 0.000 145.515 2889.180 148.245 ;
        RECT 0.000 145.465 132.745 145.515 ;
        RECT 0.000 142.805 173.225 142.855 ;
        RECT 0.000 140.075 2889.180 142.805 ;
        RECT 0.000 140.025 89.045 140.075 ;
        RECT 0.000 137.365 309.845 137.415 ;
        RECT 0.000 134.635 2889.180 137.365 ;
        RECT 0.000 134.585 47.645 134.635 ;
        RECT 0.000 131.925 90.885 131.975 ;
        RECT 0.000 129.195 2889.180 131.925 ;
        RECT 0.000 129.145 88.585 129.195 ;
        RECT 0.000 126.485 1122.665 126.535 ;
        RECT 0.000 123.755 2889.180 126.485 ;
        RECT 0.000 123.705 113.885 123.755 ;
        RECT 0.000 121.045 186.105 121.095 ;
        RECT 0.000 118.315 2889.180 121.045 ;
        RECT 0.000 118.265 141.945 118.315 ;
        RECT 0.000 115.605 279.485 115.655 ;
        RECT 0.000 112.875 2889.180 115.605 ;
        RECT 0.000 112.825 394.485 112.875 ;
        RECT 0.000 110.165 199.445 110.215 ;
        RECT 0.000 107.435 2889.180 110.165 ;
        RECT 0.000 107.385 181.505 107.435 ;
        RECT 0.000 104.725 47.645 104.775 ;
        RECT 0.000 101.995 2889.180 104.725 ;
        RECT 0.000 101.945 161.725 101.995 ;
        RECT 0.000 99.285 128.145 99.335 ;
        RECT 0.000 96.555 2889.180 99.285 ;
        RECT 0.000 96.505 703.145 96.555 ;
        RECT 0.000 93.845 201.285 93.895 ;
        RECT 0.000 91.115 2889.180 93.845 ;
        RECT 0.000 91.065 29.705 91.115 ;
        RECT 0.000 88.405 65.125 88.455 ;
        RECT 0.000 85.675 2889.180 88.405 ;
        RECT 0.000 85.625 101.005 85.675 ;
        RECT 0.000 82.965 380.685 83.015 ;
        RECT 0.000 80.235 2889.180 82.965 ;
        RECT 0.000 80.185 338.365 80.235 ;
        RECT 0.000 77.525 241.305 77.575 ;
        RECT 0.000 74.795 2889.180 77.525 ;
        RECT 0.000 74.745 123.085 74.795 ;
        RECT 0.000 72.085 33.385 72.135 ;
        RECT 0.000 69.355 2889.180 72.085 ;
        RECT 0.000 69.305 170.925 69.355 ;
        RECT 0.000 66.645 117.565 66.695 ;
        RECT 0.000 63.915 2889.180 66.645 ;
        RECT 0.000 63.865 72.025 63.915 ;
        RECT 0.000 61.205 111.585 61.255 ;
        RECT 0.000 58.475 2889.180 61.205 ;
        RECT 0.000 58.425 118.025 58.475 ;
        RECT 0.000 55.765 52.245 55.815 ;
        RECT 0.000 53.035 2889.180 55.765 ;
        RECT 0.000 52.985 57.765 53.035 ;
        RECT 0.000 50.325 167.705 50.375 ;
        RECT 0.000 47.595 2889.180 50.325 ;
        RECT 0.000 47.545 85.825 47.595 ;
        RECT 0.000 44.885 101.005 44.935 ;
        RECT 0.000 42.155 2889.180 44.885 ;
        RECT 0.000 42.105 684.745 42.155 ;
        RECT 0.000 39.445 645.185 39.495 ;
        RECT 0.000 36.715 2889.180 39.445 ;
        RECT 0.000 36.665 688.425 36.715 ;
        RECT 0.000 34.005 717.865 34.055 ;
        RECT 0.000 31.275 2889.180 34.005 ;
        RECT 0.000 31.225 794.685 31.275 ;
        RECT 0.000 28.565 808.945 28.615 ;
        RECT 0.000 25.835 2889.180 28.565 ;
        RECT 0.000 25.785 746.845 25.835 ;
        RECT 0.000 23.125 838.845 23.175 ;
        RECT 0.000 20.395 2889.180 23.125 ;
        RECT 0.000 20.345 1208.225 20.395 ;
        RECT 0.000 17.685 1176.485 17.735 ;
        RECT 0.000 14.905 2889.180 17.685 ;
        RECT 0.000 10.690 2889.180 12.295 ;
      LAYER li1 ;
        RECT 0.190 10.795 2889.765 3087.285 ;
      LAYER met1 ;
        RECT 0.190 9.900 2889.825 3087.440 ;
      LAYER met2 ;
        RECT 1.670 4.280 2887.970 3087.440 ;
        RECT 1.670 4.000 11.500 4.280 ;
        RECT 12.340 4.000 46.000 4.280 ;
        RECT 46.840 4.000 80.960 4.280 ;
        RECT 81.800 4.000 115.920 4.280 ;
        RECT 116.760 4.000 150.880 4.280 ;
        RECT 151.720 4.000 185.840 4.280 ;
        RECT 186.680 4.000 220.800 4.280 ;
        RECT 221.640 4.000 255.760 4.280 ;
        RECT 256.600 4.000 290.720 4.280 ;
        RECT 291.560 4.000 325.680 4.280 ;
        RECT 326.520 4.000 360.640 4.280 ;
        RECT 361.480 4.000 395.600 4.280 ;
        RECT 396.440 4.000 430.560 4.280 ;
        RECT 431.400 4.000 465.520 4.280 ;
        RECT 466.360 4.000 500.480 4.280 ;
        RECT 501.320 4.000 535.440 4.280 ;
        RECT 536.280 4.000 570.400 4.280 ;
        RECT 571.240 4.000 605.360 4.280 ;
        RECT 606.200 4.000 640.320 4.280 ;
        RECT 641.160 4.000 675.280 4.280 ;
        RECT 676.120 4.000 710.240 4.280 ;
        RECT 711.080 4.000 744.740 4.280 ;
        RECT 745.580 4.000 779.700 4.280 ;
        RECT 780.540 4.000 814.660 4.280 ;
        RECT 815.500 4.000 849.620 4.280 ;
        RECT 850.460 4.000 884.580 4.280 ;
        RECT 885.420 4.000 919.540 4.280 ;
        RECT 920.380 4.000 954.500 4.280 ;
        RECT 955.340 4.000 989.460 4.280 ;
        RECT 990.300 4.000 1024.420 4.280 ;
        RECT 1025.260 4.000 1059.380 4.280 ;
        RECT 1060.220 4.000 1094.340 4.280 ;
        RECT 1095.180 4.000 1129.300 4.280 ;
        RECT 1130.140 4.000 1164.260 4.280 ;
        RECT 1165.100 4.000 1199.220 4.280 ;
        RECT 1200.060 4.000 1234.180 4.280 ;
        RECT 1235.020 4.000 1269.140 4.280 ;
        RECT 1269.980 4.000 1304.100 4.280 ;
        RECT 1304.940 4.000 1339.060 4.280 ;
        RECT 1339.900 4.000 1374.020 4.280 ;
        RECT 1374.860 4.000 1408.980 4.280 ;
        RECT 1409.820 4.000 1443.940 4.280 ;
        RECT 1444.780 4.000 1478.440 4.280 ;
        RECT 1479.280 4.000 1513.400 4.280 ;
        RECT 1514.240 4.000 1548.360 4.280 ;
        RECT 1549.200 4.000 1583.320 4.280 ;
        RECT 1584.160 4.000 1618.280 4.280 ;
        RECT 1619.120 4.000 1653.240 4.280 ;
        RECT 1654.080 4.000 1688.200 4.280 ;
        RECT 1689.040 4.000 1723.160 4.280 ;
        RECT 1724.000 4.000 1758.120 4.280 ;
        RECT 1758.960 4.000 1793.080 4.280 ;
        RECT 1793.920 4.000 1828.040 4.280 ;
        RECT 1828.880 4.000 1863.000 4.280 ;
        RECT 1863.840 4.000 1897.960 4.280 ;
        RECT 1898.800 4.000 1932.920 4.280 ;
        RECT 1933.760 4.000 1967.880 4.280 ;
        RECT 1968.720 4.000 2002.840 4.280 ;
        RECT 2003.680 4.000 2037.800 4.280 ;
        RECT 2038.640 4.000 2072.760 4.280 ;
        RECT 2073.600 4.000 2107.720 4.280 ;
        RECT 2108.560 4.000 2142.680 4.280 ;
        RECT 2143.520 4.000 2177.640 4.280 ;
        RECT 2178.480 4.000 2212.140 4.280 ;
        RECT 2212.980 4.000 2247.100 4.280 ;
        RECT 2247.940 4.000 2282.060 4.280 ;
        RECT 2282.900 4.000 2317.020 4.280 ;
        RECT 2317.860 4.000 2351.980 4.280 ;
        RECT 2352.820 4.000 2386.940 4.280 ;
        RECT 2387.780 4.000 2421.900 4.280 ;
        RECT 2422.740 4.000 2456.860 4.280 ;
        RECT 2457.700 4.000 2491.820 4.280 ;
        RECT 2492.660 4.000 2526.780 4.280 ;
        RECT 2527.620 4.000 2561.740 4.280 ;
        RECT 2562.580 4.000 2596.700 4.280 ;
        RECT 2597.540 4.000 2631.660 4.280 ;
        RECT 2632.500 4.000 2666.620 4.280 ;
        RECT 2667.460 4.000 2701.580 4.280 ;
        RECT 2702.420 4.000 2736.540 4.280 ;
        RECT 2737.380 4.000 2771.500 4.280 ;
        RECT 2772.340 4.000 2806.460 4.280 ;
        RECT 2807.300 4.000 2841.420 4.280 ;
        RECT 2842.260 4.000 2876.380 4.280 ;
        RECT 2877.220 4.000 2887.970 4.280 ;
      LAYER met3 ;
        RECT 4.855 10.715 2887.085 3087.365 ;
      LAYER met4 ;
        RECT 17.965 13.095 92.110 3056.425 ;
        RECT 94.510 13.095 168.910 3056.425 ;
        RECT 171.310 13.095 245.710 3056.425 ;
        RECT 248.110 13.095 322.510 3056.425 ;
        RECT 324.910 13.095 399.310 3056.425 ;
        RECT 401.710 13.095 476.110 3056.425 ;
        RECT 478.510 13.095 552.910 3056.425 ;
        RECT 555.310 13.095 629.710 3056.425 ;
        RECT 632.110 13.095 706.510 3056.425 ;
        RECT 708.910 13.095 783.310 3056.425 ;
        RECT 785.710 13.095 860.110 3056.425 ;
        RECT 862.510 13.095 936.910 3056.425 ;
        RECT 939.310 13.095 1013.710 3056.425 ;
        RECT 1016.110 13.095 1090.510 3056.425 ;
        RECT 1092.910 13.095 1167.310 3056.425 ;
        RECT 1169.710 13.095 1244.110 3056.425 ;
        RECT 1246.510 13.095 1320.910 3056.425 ;
        RECT 1323.310 13.095 1397.710 3056.425 ;
        RECT 1400.110 13.095 1474.510 3056.425 ;
        RECT 1476.910 13.095 1551.310 3056.425 ;
        RECT 1553.710 13.095 1628.110 3056.425 ;
        RECT 1630.510 13.095 1704.910 3056.425 ;
        RECT 1707.310 13.095 1781.710 3056.425 ;
        RECT 1784.110 13.095 1858.510 3056.425 ;
        RECT 1860.910 13.095 1935.310 3056.425 ;
        RECT 1937.710 13.095 2012.110 3056.425 ;
        RECT 2014.510 13.095 2088.910 3056.425 ;
        RECT 2091.310 13.095 2165.710 3056.425 ;
        RECT 2168.110 13.095 2242.510 3056.425 ;
        RECT 2244.910 13.095 2319.310 3056.425 ;
        RECT 2321.710 13.095 2396.110 3056.425 ;
        RECT 2398.510 13.095 2472.910 3056.425 ;
        RECT 2475.310 13.095 2549.710 3056.425 ;
        RECT 2552.110 13.095 2626.510 3056.425 ;
        RECT 2628.910 13.095 2703.310 3056.425 ;
        RECT 2705.710 13.095 2780.110 3056.425 ;
        RECT 2782.510 13.095 2806.815 3056.425 ;
  END
END RAM_6Kx32
END LIBRARY

