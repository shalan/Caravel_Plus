VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3519.700 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3519.700 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3519.700 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3519.700 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3519.700 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3519.700 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3519.700 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3519.700 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3519.700 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 0.300 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 0.300 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 0.300 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 0.300 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 0.300 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 0.300 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 0.300 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2433.460 2924.800 2434.660 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2903.340 2924.800 2904.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3519.700 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3519.700 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3519.700 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3519.700 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3519.700 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3519.700 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3519.700 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3519.700 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3519.700 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3410.620 0.300 3411.820 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 0.300 3124.860 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2836.020 0.300 2837.220 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 0.300 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 0.300 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1974.460 0.300 1975.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 0.300 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 0.300 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 0.300 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 0.300 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 0.300 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 0.300 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 0.300 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 0.300 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1964.260 2924.800 1965.460 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2198.860 2924.800 2200.060 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3519.700 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3519.700 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3519.700 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3519.700 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3519.700 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3519.700 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3519.700 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3519.700 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3519.700 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 0.300 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 0.300 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 0.300 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 0.300 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 0.300 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 0.300 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 0.300 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 0.300 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 0.300 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 0.300 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 0.300 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 0.300 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 0.300 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 0.300 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3519.700 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3519.700 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3519.700 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3519.700 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3519.700 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3519.700 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3519.700 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3519.700 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3519.700 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.220 0.300 3340.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 0.300 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 0.300 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2476.980 0.300 2478.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 0.300 2190.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 0.300 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 0.300 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 0.300 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 0.300 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 0.300 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 0.300 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 0.300 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 0.300 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 0.300 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 0.300 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 0.300 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 0.300 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 0.300 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 0.300 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 0.300 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 0.300 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 0.300 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 0.300 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 0.300 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 0.300 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 0.300 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 0.300 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 0.300 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 0.300 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 0.300 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 0.300 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 0.300 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 0.300 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 0.300 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 0.300 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 0.300 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 0.300 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 0.300 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 0.300 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 0.300 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 0.300 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 0.300 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 0.300 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 0.300 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 0.300 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 0.300 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 0.300 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 0.300 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 0.300 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 0.300 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 0.300 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 0.300 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 0.300 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 0.300 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 0.300 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 0.300 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 0.300 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 0.300 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 0.300 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 0.300 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 0.300 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 0.300 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 0.300 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 0.300 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 0.300 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 0.300 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 0.300 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 0.300 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 0.300 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 0.300 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 0.300 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 0.300 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 0.300 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 0.300 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 0.300 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 0.300 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 0.300 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 0.300 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 0.300 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 0.300 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 0.300 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 0.300 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 0.300 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 0.300 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 0.300 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 0.300 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 0.300 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 0.300 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 0.300 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 0.300 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 0.300 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 0.300 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 0.300 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 0.300 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 0.300 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 0.300 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 0.300 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 0.300 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 0.300 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 0.300 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 0.300 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 0.300 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 0.300 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 0.300 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 0.300 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 0.300 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 0.300 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 0.300 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 0.300 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 0.300 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 0.300 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 0.300 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 0.300 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 0.300 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 0.300 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 0.300 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 0.300 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 0.300 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 0.300 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 0.300 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 0.300 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 0.300 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 0.300 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 0.300 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 0.300 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 0.300 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 0.300 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 0.300 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 0.300 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 0.300 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 0.300 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 0.300 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 0.300 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 0.300 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 0.300 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 0.300 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 0.300 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 0.300 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 0.300 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 0.300 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 0.300 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 0.300 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 0.300 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 0.300 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 0.300 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 0.300 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 0.300 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 0.300 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 0.300 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 0.300 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 0.300 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 0.300 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 0.300 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 0.300 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 0.300 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 0.300 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 0.300 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 0.300 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 0.300 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 0.300 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 0.300 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 0.300 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 0.300 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 0.300 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 0.300 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 0.300 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 0.300 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 0.300 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 0.300 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 0.300 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 0.300 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 0.300 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 0.300 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 0.300 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 0.300 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 0.300 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 0.300 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 0.300 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 0.300 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 0.300 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 0.300 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 0.300 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 0.300 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 0.300 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 0.300 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 0.300 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 0.300 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 0.300 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 0.300 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 0.300 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 0.300 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 0.300 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 0.300 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 0.300 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 0.300 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 0.300 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 0.300 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 0.300 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 0.300 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 0.300 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 0.300 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 0.300 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 0.300 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 0.300 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 0.300 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 0.300 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 0.300 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 0.300 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 0.300 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 0.300 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 0.300 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 0.300 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 0.300 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 0.300 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 0.300 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 0.300 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 0.300 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 0.300 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 0.300 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 0.300 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 0.300 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 0.300 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 0.300 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 0.300 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 0.300 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 0.300 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 0.300 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 0.300 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 0.300 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 0.300 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 0.300 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 0.300 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 0.300 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 0.300 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 0.300 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 0.300 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 0.300 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 0.300 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 0.300 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 0.300 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 0.300 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 0.300 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 0.300 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 0.300 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 0.300 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 0.300 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 0.300 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 0.300 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 0.300 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 0.300 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 0.300 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 0.300 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 0.300 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 0.300 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 0.300 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 0.300 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 0.300 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 0.300 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 0.300 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 0.300 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 0.300 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 0.300 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 0.300 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 0.300 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 0.300 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 0.300 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 0.300 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 0.300 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 0.300 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 0.300 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 0.300 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 0.300 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 0.300 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 0.300 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 0.300 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 0.300 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 0.300 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 0.300 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 0.300 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 0.300 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 0.300 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 0.300 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 0.300 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 0.300 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 0.300 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 0.300 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 0.300 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 0.300 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 0.300 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 0.300 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 0.300 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 0.300 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 0.300 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 0.300 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 0.300 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 0.300 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 0.300 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 0.300 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 0.300 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 0.300 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 0.300 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 0.300 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 0.300 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 0.300 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 0.300 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 0.300 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 0.300 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 0.300 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 0.300 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 0.300 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 0.300 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 0.300 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 0.300 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 0.300 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 0.300 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 0.300 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 0.300 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 0.300 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 0.300 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 0.300 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 0.300 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 0.300 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 0.300 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 0.300 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 0.300 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 0.300 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 0.300 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 0.300 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 0.300 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 0.300 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 0.300 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 0.300 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 0.300 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 0.300 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 0.300 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 0.300 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 0.300 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 0.300 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 0.300 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 0.300 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 0.300 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 0.300 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 0.300 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 0.300 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 0.300 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 0.300 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 0.300 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 0.300 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 0.300 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 0.300 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 0.300 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 0.300 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 0.300 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 0.300 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 0.300 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 0.300 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 0.300 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 0.300 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 0.300 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 0.300 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 0.300 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 0.300 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 0.300 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 0.300 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 0.300 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 0.300 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 0.300 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 0.300 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 0.300 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 0.300 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 0.300 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 0.300 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 0.300 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 0.300 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 0.300 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 0.300 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 0.300 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 0.300 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 0.300 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 0.300 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 0.300 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 0.300 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 0.300 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 0.300 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 0.300 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 0.300 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 0.300 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 0.300 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 0.300 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 0.300 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 0.300 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 0.300 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 0.300 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 0.300 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 0.300 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 0.300 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 0.300 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 0.300 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 0.300 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 0.300 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 0.300 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 0.300 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 0.300 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 0.300 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 0.300 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 0.300 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 0.300 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 0.300 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 0.300 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 0.300 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 0.300 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 0.300 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 0.300 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 0.300 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 0.300 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 0.300 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 0.300 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 0.300 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 0.300 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 0.300 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 0.300 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 0.300 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 0.300 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 0.300 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 0.300 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 0.300 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 0.300 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 0.300 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 0.300 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 0.300 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 0.300 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 0.300 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 0.300 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 0.300 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 0.300 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 0.300 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 0.300 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 0.300 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 0.300 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 0.300 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 0.300 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 0.300 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 0.300 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 0.300 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 0.300 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 0.300 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 0.300 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 0.300 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 0.300 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 0.300 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 0.300 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 0.300 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 0.300 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 0.300 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 0.300 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 0.300 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 0.300 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 0.300 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 0.300 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 0.300 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 0.300 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 0.300 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 0.300 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 0.300 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 0.300 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 0.300 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 0.300 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 0.300 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 0.300 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 0.300 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 0.300 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 0.300 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 0.300 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 0.300 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 0.300 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 0.300 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 0.300 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 0.300 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 0.300 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 0.300 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 0.300 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 0.300 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 0.300 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 0.300 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 0.300 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 0.300 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 0.300 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 0.300 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 0.300 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 0.300 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 0.300 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 0.300 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 0.300 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 0.300 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 0.300 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 0.300 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 0.300 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 0.300 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 0.300 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 0.300 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 0.300 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 0.300 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 0.300 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 0.300 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 0.300 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 3519.700 7.020 3528.900 ;
        RECT 184.020 3519.700 187.020 3528.900 ;
        RECT 364.020 3519.700 367.020 3528.900 ;
        RECT 544.020 3519.700 547.020 3528.900 ;
        RECT 724.020 3519.700 727.020 3528.900 ;
        RECT 904.020 3519.700 907.020 3528.900 ;
        RECT 1084.020 3519.700 1087.020 3528.900 ;
        RECT 1264.020 3519.700 1267.020 3528.900 ;
        RECT 1444.020 3519.700 1447.020 3528.900 ;
        RECT 1624.020 3519.700 1627.020 3528.900 ;
        RECT 1804.020 3519.700 1807.020 3528.900 ;
        RECT 1984.020 3519.700 1987.020 3528.900 ;
        RECT 2164.020 3519.700 2167.020 3528.900 ;
        RECT 2344.020 3519.700 2347.020 3528.900 ;
        RECT 2524.020 3519.700 2527.020 3528.900 ;
        RECT 2704.020 3519.700 2707.020 3528.900 ;
        RECT 2884.020 3519.700 2887.020 3528.900 ;
        RECT 4.020 -9.220 7.020 0.300 ;
        RECT 184.020 -9.220 187.020 0.300 ;
        RECT 364.020 -9.220 367.020 0.300 ;
        RECT 544.020 -9.220 547.020 0.300 ;
        RECT 724.020 -9.220 727.020 0.300 ;
        RECT 904.020 -9.220 907.020 0.300 ;
        RECT 1084.020 -9.220 1087.020 0.300 ;
        RECT 1264.020 -9.220 1267.020 0.300 ;
        RECT 1444.020 -9.220 1447.020 0.300 ;
        RECT 1624.020 -9.220 1627.020 0.300 ;
        RECT 1804.020 -9.220 1807.020 0.300 ;
        RECT 1984.020 -9.220 1987.020 0.300 ;
        RECT 2164.020 -9.220 2167.020 0.300 ;
        RECT 2344.020 -9.220 2347.020 0.300 ;
        RECT 2524.020 -9.220 2527.020 0.300 ;
        RECT 2704.020 -9.220 2707.020 0.300 ;
        RECT 2884.020 -9.220 2887.020 0.300 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT -9.070 3430.850 -7.890 3432.030 ;
        RECT -9.070 3429.250 -7.890 3430.430 ;
        RECT -9.070 3250.850 -7.890 3252.030 ;
        RECT -9.070 3249.250 -7.890 3250.430 ;
        RECT -9.070 3070.850 -7.890 3072.030 ;
        RECT -9.070 3069.250 -7.890 3070.430 ;
        RECT -9.070 2890.850 -7.890 2892.030 ;
        RECT -9.070 2889.250 -7.890 2890.430 ;
        RECT -9.070 2710.850 -7.890 2712.030 ;
        RECT -9.070 2709.250 -7.890 2710.430 ;
        RECT -9.070 2530.850 -7.890 2532.030 ;
        RECT -9.070 2529.250 -7.890 2530.430 ;
        RECT -9.070 2350.850 -7.890 2352.030 ;
        RECT -9.070 2349.250 -7.890 2350.430 ;
        RECT -9.070 2170.850 -7.890 2172.030 ;
        RECT -9.070 2169.250 -7.890 2170.430 ;
        RECT -9.070 1990.850 -7.890 1992.030 ;
        RECT -9.070 1989.250 -7.890 1990.430 ;
        RECT -9.070 1810.850 -7.890 1812.030 ;
        RECT -9.070 1809.250 -7.890 1810.430 ;
        RECT -9.070 1630.850 -7.890 1632.030 ;
        RECT -9.070 1629.250 -7.890 1630.430 ;
        RECT -9.070 1450.850 -7.890 1452.030 ;
        RECT -9.070 1449.250 -7.890 1450.430 ;
        RECT -9.070 1270.850 -7.890 1272.030 ;
        RECT -9.070 1269.250 -7.890 1270.430 ;
        RECT -9.070 1090.850 -7.890 1092.030 ;
        RECT -9.070 1089.250 -7.890 1090.430 ;
        RECT -9.070 910.850 -7.890 912.030 ;
        RECT -9.070 909.250 -7.890 910.430 ;
        RECT -9.070 730.850 -7.890 732.030 ;
        RECT -9.070 729.250 -7.890 730.430 ;
        RECT -9.070 550.850 -7.890 552.030 ;
        RECT -9.070 549.250 -7.890 550.430 ;
        RECT -9.070 370.850 -7.890 372.030 ;
        RECT -9.070 369.250 -7.890 370.430 ;
        RECT -9.070 190.850 -7.890 192.030 ;
        RECT -9.070 189.250 -7.890 190.430 ;
        RECT -9.070 10.850 -7.890 12.030 ;
        RECT -9.070 9.250 -7.890 10.430 ;
        RECT 2927.510 3430.850 2928.690 3432.030 ;
        RECT 2927.510 3429.250 2928.690 3430.430 ;
        RECT 2927.510 3250.850 2928.690 3252.030 ;
        RECT 2927.510 3249.250 2928.690 3250.430 ;
        RECT 2927.510 3070.850 2928.690 3072.030 ;
        RECT 2927.510 3069.250 2928.690 3070.430 ;
        RECT 2927.510 2890.850 2928.690 2892.030 ;
        RECT 2927.510 2889.250 2928.690 2890.430 ;
        RECT 2927.510 2710.850 2928.690 2712.030 ;
        RECT 2927.510 2709.250 2928.690 2710.430 ;
        RECT 2927.510 2530.850 2928.690 2532.030 ;
        RECT 2927.510 2529.250 2928.690 2530.430 ;
        RECT 2927.510 2350.850 2928.690 2352.030 ;
        RECT 2927.510 2349.250 2928.690 2350.430 ;
        RECT 2927.510 2170.850 2928.690 2172.030 ;
        RECT 2927.510 2169.250 2928.690 2170.430 ;
        RECT 2927.510 1990.850 2928.690 1992.030 ;
        RECT 2927.510 1989.250 2928.690 1990.430 ;
        RECT 2927.510 1810.850 2928.690 1812.030 ;
        RECT 2927.510 1809.250 2928.690 1810.430 ;
        RECT 2927.510 1630.850 2928.690 1632.030 ;
        RECT 2927.510 1629.250 2928.690 1630.430 ;
        RECT 2927.510 1450.850 2928.690 1452.030 ;
        RECT 2927.510 1449.250 2928.690 1450.430 ;
        RECT 2927.510 1270.850 2928.690 1272.030 ;
        RECT 2927.510 1269.250 2928.690 1270.430 ;
        RECT 2927.510 1090.850 2928.690 1092.030 ;
        RECT 2927.510 1089.250 2928.690 1090.430 ;
        RECT 2927.510 910.850 2928.690 912.030 ;
        RECT 2927.510 909.250 2928.690 910.430 ;
        RECT 2927.510 730.850 2928.690 732.030 ;
        RECT 2927.510 729.250 2928.690 730.430 ;
        RECT 2927.510 550.850 2928.690 552.030 ;
        RECT 2927.510 549.250 2928.690 550.430 ;
        RECT 2927.510 370.850 2928.690 372.030 ;
        RECT 2927.510 369.250 2928.690 370.430 ;
        RECT 2927.510 190.850 2928.690 192.030 ;
        RECT 2927.510 189.250 2928.690 190.430 ;
        RECT 2927.510 10.850 2928.690 12.030 ;
        RECT 2927.510 9.250 2928.690 10.430 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.140 -6.980 3432.150 ;
        RECT 2926.600 3432.140 2929.600 3432.150 ;
        RECT -14.580 3429.140 0.300 3432.140 ;
        RECT 2919.700 3429.140 2934.200 3432.140 ;
        RECT -9.980 3429.130 -6.980 3429.140 ;
        RECT 2926.600 3429.130 2929.600 3429.140 ;
        RECT -9.980 3252.140 -6.980 3252.150 ;
        RECT 2926.600 3252.140 2929.600 3252.150 ;
        RECT -14.580 3249.140 0.300 3252.140 ;
        RECT 2919.700 3249.140 2934.200 3252.140 ;
        RECT -9.980 3249.130 -6.980 3249.140 ;
        RECT 2926.600 3249.130 2929.600 3249.140 ;
        RECT -9.980 3072.140 -6.980 3072.150 ;
        RECT 2926.600 3072.140 2929.600 3072.150 ;
        RECT -14.580 3069.140 0.300 3072.140 ;
        RECT 2919.700 3069.140 2934.200 3072.140 ;
        RECT -9.980 3069.130 -6.980 3069.140 ;
        RECT 2926.600 3069.130 2929.600 3069.140 ;
        RECT -9.980 2892.140 -6.980 2892.150 ;
        RECT 2926.600 2892.140 2929.600 2892.150 ;
        RECT -14.580 2889.140 0.300 2892.140 ;
        RECT 2919.700 2889.140 2934.200 2892.140 ;
        RECT -9.980 2889.130 -6.980 2889.140 ;
        RECT 2926.600 2889.130 2929.600 2889.140 ;
        RECT -9.980 2712.140 -6.980 2712.150 ;
        RECT 2926.600 2712.140 2929.600 2712.150 ;
        RECT -14.580 2709.140 0.300 2712.140 ;
        RECT 2919.700 2709.140 2934.200 2712.140 ;
        RECT -9.980 2709.130 -6.980 2709.140 ;
        RECT 2926.600 2709.130 2929.600 2709.140 ;
        RECT -9.980 2532.140 -6.980 2532.150 ;
        RECT 2926.600 2532.140 2929.600 2532.150 ;
        RECT -14.580 2529.140 0.300 2532.140 ;
        RECT 2919.700 2529.140 2934.200 2532.140 ;
        RECT -9.980 2529.130 -6.980 2529.140 ;
        RECT 2926.600 2529.130 2929.600 2529.140 ;
        RECT -9.980 2352.140 -6.980 2352.150 ;
        RECT 2926.600 2352.140 2929.600 2352.150 ;
        RECT -14.580 2349.140 0.300 2352.140 ;
        RECT 2919.700 2349.140 2934.200 2352.140 ;
        RECT -9.980 2349.130 -6.980 2349.140 ;
        RECT 2926.600 2349.130 2929.600 2349.140 ;
        RECT -9.980 2172.140 -6.980 2172.150 ;
        RECT 2926.600 2172.140 2929.600 2172.150 ;
        RECT -14.580 2169.140 0.300 2172.140 ;
        RECT 2919.700 2169.140 2934.200 2172.140 ;
        RECT -9.980 2169.130 -6.980 2169.140 ;
        RECT 2926.600 2169.130 2929.600 2169.140 ;
        RECT -9.980 1992.140 -6.980 1992.150 ;
        RECT 2926.600 1992.140 2929.600 1992.150 ;
        RECT -14.580 1989.140 0.300 1992.140 ;
        RECT 2919.700 1989.140 2934.200 1992.140 ;
        RECT -9.980 1989.130 -6.980 1989.140 ;
        RECT 2926.600 1989.130 2929.600 1989.140 ;
        RECT -9.980 1812.140 -6.980 1812.150 ;
        RECT 2926.600 1812.140 2929.600 1812.150 ;
        RECT -14.580 1809.140 0.300 1812.140 ;
        RECT 2919.700 1809.140 2934.200 1812.140 ;
        RECT -9.980 1809.130 -6.980 1809.140 ;
        RECT 2926.600 1809.130 2929.600 1809.140 ;
        RECT -9.980 1632.140 -6.980 1632.150 ;
        RECT 2926.600 1632.140 2929.600 1632.150 ;
        RECT -14.580 1629.140 0.300 1632.140 ;
        RECT 2919.700 1629.140 2934.200 1632.140 ;
        RECT -9.980 1629.130 -6.980 1629.140 ;
        RECT 2926.600 1629.130 2929.600 1629.140 ;
        RECT -9.980 1452.140 -6.980 1452.150 ;
        RECT 2926.600 1452.140 2929.600 1452.150 ;
        RECT -14.580 1449.140 0.300 1452.140 ;
        RECT 2919.700 1449.140 2934.200 1452.140 ;
        RECT -9.980 1449.130 -6.980 1449.140 ;
        RECT 2926.600 1449.130 2929.600 1449.140 ;
        RECT -9.980 1272.140 -6.980 1272.150 ;
        RECT 2926.600 1272.140 2929.600 1272.150 ;
        RECT -14.580 1269.140 0.300 1272.140 ;
        RECT 2919.700 1269.140 2934.200 1272.140 ;
        RECT -9.980 1269.130 -6.980 1269.140 ;
        RECT 2926.600 1269.130 2929.600 1269.140 ;
        RECT -9.980 1092.140 -6.980 1092.150 ;
        RECT 2926.600 1092.140 2929.600 1092.150 ;
        RECT -14.580 1089.140 0.300 1092.140 ;
        RECT 2919.700 1089.140 2934.200 1092.140 ;
        RECT -9.980 1089.130 -6.980 1089.140 ;
        RECT 2926.600 1089.130 2929.600 1089.140 ;
        RECT -9.980 912.140 -6.980 912.150 ;
        RECT 2926.600 912.140 2929.600 912.150 ;
        RECT -14.580 909.140 0.300 912.140 ;
        RECT 2919.700 909.140 2934.200 912.140 ;
        RECT -9.980 909.130 -6.980 909.140 ;
        RECT 2926.600 909.130 2929.600 909.140 ;
        RECT -9.980 732.140 -6.980 732.150 ;
        RECT 2926.600 732.140 2929.600 732.150 ;
        RECT -14.580 729.140 0.300 732.140 ;
        RECT 2919.700 729.140 2934.200 732.140 ;
        RECT -9.980 729.130 -6.980 729.140 ;
        RECT 2926.600 729.130 2929.600 729.140 ;
        RECT -9.980 552.140 -6.980 552.150 ;
        RECT 2926.600 552.140 2929.600 552.150 ;
        RECT -14.580 549.140 0.300 552.140 ;
        RECT 2919.700 549.140 2934.200 552.140 ;
        RECT -9.980 549.130 -6.980 549.140 ;
        RECT 2926.600 549.130 2929.600 549.140 ;
        RECT -9.980 372.140 -6.980 372.150 ;
        RECT 2926.600 372.140 2929.600 372.150 ;
        RECT -14.580 369.140 0.300 372.140 ;
        RECT 2919.700 369.140 2934.200 372.140 ;
        RECT -9.980 369.130 -6.980 369.140 ;
        RECT 2926.600 369.130 2929.600 369.140 ;
        RECT -9.980 192.140 -6.980 192.150 ;
        RECT 2926.600 192.140 2929.600 192.150 ;
        RECT -14.580 189.140 0.300 192.140 ;
        RECT 2919.700 189.140 2934.200 192.140 ;
        RECT -9.980 189.130 -6.980 189.140 ;
        RECT 2926.600 189.130 2929.600 189.140 ;
        RECT -9.980 12.140 -6.980 12.150 ;
        RECT 2926.600 12.140 2929.600 12.150 ;
        RECT -14.580 9.140 0.300 12.140 ;
        RECT 2919.700 9.140 2934.200 12.140 ;
        RECT -9.980 9.130 -6.980 9.140 ;
        RECT 2926.600 9.130 2929.600 9.140 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 3519.700 97.020 3528.900 ;
        RECT 274.020 3519.700 277.020 3528.900 ;
        RECT 454.020 3519.700 457.020 3528.900 ;
        RECT 634.020 3519.700 637.020 3528.900 ;
        RECT 814.020 3519.700 817.020 3528.900 ;
        RECT 994.020 3519.700 997.020 3528.900 ;
        RECT 1174.020 3519.700 1177.020 3528.900 ;
        RECT 1354.020 3519.700 1357.020 3528.900 ;
        RECT 1534.020 3519.700 1537.020 3528.900 ;
        RECT 1714.020 3519.700 1717.020 3528.900 ;
        RECT 1894.020 3519.700 1897.020 3528.900 ;
        RECT 2074.020 3519.700 2077.020 3528.900 ;
        RECT 2254.020 3519.700 2257.020 3528.900 ;
        RECT 2434.020 3519.700 2437.020 3528.900 ;
        RECT 2614.020 3519.700 2617.020 3528.900 ;
        RECT 2794.020 3519.700 2797.020 3528.900 ;
        RECT 94.020 -9.220 97.020 0.300 ;
        RECT 274.020 -9.220 277.020 0.300 ;
        RECT 454.020 -9.220 457.020 0.300 ;
        RECT 634.020 -9.220 637.020 0.300 ;
        RECT 814.020 -9.220 817.020 0.300 ;
        RECT 994.020 -9.220 997.020 0.300 ;
        RECT 1174.020 -9.220 1177.020 0.300 ;
        RECT 1354.020 -9.220 1357.020 0.300 ;
        RECT 1534.020 -9.220 1537.020 0.300 ;
        RECT 1714.020 -9.220 1717.020 0.300 ;
        RECT 1894.020 -9.220 1897.020 0.300 ;
        RECT 2074.020 -9.220 2077.020 0.300 ;
        RECT 2254.020 -9.220 2257.020 0.300 ;
        RECT 2434.020 -9.220 2437.020 0.300 ;
        RECT 2614.020 -9.220 2617.020 0.300 ;
        RECT 2794.020 -9.220 2797.020 0.300 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT -13.670 3340.850 -12.490 3342.030 ;
        RECT -13.670 3339.250 -12.490 3340.430 ;
        RECT -13.670 3160.850 -12.490 3162.030 ;
        RECT -13.670 3159.250 -12.490 3160.430 ;
        RECT -13.670 2980.850 -12.490 2982.030 ;
        RECT -13.670 2979.250 -12.490 2980.430 ;
        RECT -13.670 2800.850 -12.490 2802.030 ;
        RECT -13.670 2799.250 -12.490 2800.430 ;
        RECT -13.670 2620.850 -12.490 2622.030 ;
        RECT -13.670 2619.250 -12.490 2620.430 ;
        RECT -13.670 2440.850 -12.490 2442.030 ;
        RECT -13.670 2439.250 -12.490 2440.430 ;
        RECT -13.670 2260.850 -12.490 2262.030 ;
        RECT -13.670 2259.250 -12.490 2260.430 ;
        RECT -13.670 2080.850 -12.490 2082.030 ;
        RECT -13.670 2079.250 -12.490 2080.430 ;
        RECT -13.670 1900.850 -12.490 1902.030 ;
        RECT -13.670 1899.250 -12.490 1900.430 ;
        RECT -13.670 1720.850 -12.490 1722.030 ;
        RECT -13.670 1719.250 -12.490 1720.430 ;
        RECT -13.670 1540.850 -12.490 1542.030 ;
        RECT -13.670 1539.250 -12.490 1540.430 ;
        RECT -13.670 1360.850 -12.490 1362.030 ;
        RECT -13.670 1359.250 -12.490 1360.430 ;
        RECT -13.670 1180.850 -12.490 1182.030 ;
        RECT -13.670 1179.250 -12.490 1180.430 ;
        RECT -13.670 1000.850 -12.490 1002.030 ;
        RECT -13.670 999.250 -12.490 1000.430 ;
        RECT -13.670 820.850 -12.490 822.030 ;
        RECT -13.670 819.250 -12.490 820.430 ;
        RECT -13.670 640.850 -12.490 642.030 ;
        RECT -13.670 639.250 -12.490 640.430 ;
        RECT -13.670 460.850 -12.490 462.030 ;
        RECT -13.670 459.250 -12.490 460.430 ;
        RECT -13.670 280.850 -12.490 282.030 ;
        RECT -13.670 279.250 -12.490 280.430 ;
        RECT -13.670 100.850 -12.490 102.030 ;
        RECT -13.670 99.250 -12.490 100.430 ;
        RECT 2932.110 3340.850 2933.290 3342.030 ;
        RECT 2932.110 3339.250 2933.290 3340.430 ;
        RECT 2932.110 3160.850 2933.290 3162.030 ;
        RECT 2932.110 3159.250 2933.290 3160.430 ;
        RECT 2932.110 2980.850 2933.290 2982.030 ;
        RECT 2932.110 2979.250 2933.290 2980.430 ;
        RECT 2932.110 2800.850 2933.290 2802.030 ;
        RECT 2932.110 2799.250 2933.290 2800.430 ;
        RECT 2932.110 2620.850 2933.290 2622.030 ;
        RECT 2932.110 2619.250 2933.290 2620.430 ;
        RECT 2932.110 2440.850 2933.290 2442.030 ;
        RECT 2932.110 2439.250 2933.290 2440.430 ;
        RECT 2932.110 2260.850 2933.290 2262.030 ;
        RECT 2932.110 2259.250 2933.290 2260.430 ;
        RECT 2932.110 2080.850 2933.290 2082.030 ;
        RECT 2932.110 2079.250 2933.290 2080.430 ;
        RECT 2932.110 1900.850 2933.290 1902.030 ;
        RECT 2932.110 1899.250 2933.290 1900.430 ;
        RECT 2932.110 1720.850 2933.290 1722.030 ;
        RECT 2932.110 1719.250 2933.290 1720.430 ;
        RECT 2932.110 1540.850 2933.290 1542.030 ;
        RECT 2932.110 1539.250 2933.290 1540.430 ;
        RECT 2932.110 1360.850 2933.290 1362.030 ;
        RECT 2932.110 1359.250 2933.290 1360.430 ;
        RECT 2932.110 1180.850 2933.290 1182.030 ;
        RECT 2932.110 1179.250 2933.290 1180.430 ;
        RECT 2932.110 1000.850 2933.290 1002.030 ;
        RECT 2932.110 999.250 2933.290 1000.430 ;
        RECT 2932.110 820.850 2933.290 822.030 ;
        RECT 2932.110 819.250 2933.290 820.430 ;
        RECT 2932.110 640.850 2933.290 642.030 ;
        RECT 2932.110 639.250 2933.290 640.430 ;
        RECT 2932.110 460.850 2933.290 462.030 ;
        RECT 2932.110 459.250 2933.290 460.430 ;
        RECT 2932.110 280.850 2933.290 282.030 ;
        RECT 2932.110 279.250 2933.290 280.430 ;
        RECT 2932.110 100.850 2933.290 102.030 ;
        RECT 2932.110 99.250 2933.290 100.430 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.140 -11.580 3342.150 ;
        RECT 2931.200 3342.140 2934.200 3342.150 ;
        RECT -14.580 3339.140 0.300 3342.140 ;
        RECT 2919.700 3339.140 2934.200 3342.140 ;
        RECT -14.580 3339.130 -11.580 3339.140 ;
        RECT 2931.200 3339.130 2934.200 3339.140 ;
        RECT -14.580 3162.140 -11.580 3162.150 ;
        RECT 2931.200 3162.140 2934.200 3162.150 ;
        RECT -14.580 3159.140 0.300 3162.140 ;
        RECT 2919.700 3159.140 2934.200 3162.140 ;
        RECT -14.580 3159.130 -11.580 3159.140 ;
        RECT 2931.200 3159.130 2934.200 3159.140 ;
        RECT -14.580 2982.140 -11.580 2982.150 ;
        RECT 2931.200 2982.140 2934.200 2982.150 ;
        RECT -14.580 2979.140 0.300 2982.140 ;
        RECT 2919.700 2979.140 2934.200 2982.140 ;
        RECT -14.580 2979.130 -11.580 2979.140 ;
        RECT 2931.200 2979.130 2934.200 2979.140 ;
        RECT -14.580 2802.140 -11.580 2802.150 ;
        RECT 2931.200 2802.140 2934.200 2802.150 ;
        RECT -14.580 2799.140 0.300 2802.140 ;
        RECT 2919.700 2799.140 2934.200 2802.140 ;
        RECT -14.580 2799.130 -11.580 2799.140 ;
        RECT 2931.200 2799.130 2934.200 2799.140 ;
        RECT -14.580 2622.140 -11.580 2622.150 ;
        RECT 2931.200 2622.140 2934.200 2622.150 ;
        RECT -14.580 2619.140 0.300 2622.140 ;
        RECT 2919.700 2619.140 2934.200 2622.140 ;
        RECT -14.580 2619.130 -11.580 2619.140 ;
        RECT 2931.200 2619.130 2934.200 2619.140 ;
        RECT -14.580 2442.140 -11.580 2442.150 ;
        RECT 2931.200 2442.140 2934.200 2442.150 ;
        RECT -14.580 2439.140 0.300 2442.140 ;
        RECT 2919.700 2439.140 2934.200 2442.140 ;
        RECT -14.580 2439.130 -11.580 2439.140 ;
        RECT 2931.200 2439.130 2934.200 2439.140 ;
        RECT -14.580 2262.140 -11.580 2262.150 ;
        RECT 2931.200 2262.140 2934.200 2262.150 ;
        RECT -14.580 2259.140 0.300 2262.140 ;
        RECT 2919.700 2259.140 2934.200 2262.140 ;
        RECT -14.580 2259.130 -11.580 2259.140 ;
        RECT 2931.200 2259.130 2934.200 2259.140 ;
        RECT -14.580 2082.140 -11.580 2082.150 ;
        RECT 2931.200 2082.140 2934.200 2082.150 ;
        RECT -14.580 2079.140 0.300 2082.140 ;
        RECT 2919.700 2079.140 2934.200 2082.140 ;
        RECT -14.580 2079.130 -11.580 2079.140 ;
        RECT 2931.200 2079.130 2934.200 2079.140 ;
        RECT -14.580 1902.140 -11.580 1902.150 ;
        RECT 2931.200 1902.140 2934.200 1902.150 ;
        RECT -14.580 1899.140 0.300 1902.140 ;
        RECT 2919.700 1899.140 2934.200 1902.140 ;
        RECT -14.580 1899.130 -11.580 1899.140 ;
        RECT 2931.200 1899.130 2934.200 1899.140 ;
        RECT -14.580 1722.140 -11.580 1722.150 ;
        RECT 2931.200 1722.140 2934.200 1722.150 ;
        RECT -14.580 1719.140 0.300 1722.140 ;
        RECT 2919.700 1719.140 2934.200 1722.140 ;
        RECT -14.580 1719.130 -11.580 1719.140 ;
        RECT 2931.200 1719.130 2934.200 1719.140 ;
        RECT -14.580 1542.140 -11.580 1542.150 ;
        RECT 2931.200 1542.140 2934.200 1542.150 ;
        RECT -14.580 1539.140 0.300 1542.140 ;
        RECT 2919.700 1539.140 2934.200 1542.140 ;
        RECT -14.580 1539.130 -11.580 1539.140 ;
        RECT 2931.200 1539.130 2934.200 1539.140 ;
        RECT -14.580 1362.140 -11.580 1362.150 ;
        RECT 2931.200 1362.140 2934.200 1362.150 ;
        RECT -14.580 1359.140 0.300 1362.140 ;
        RECT 2919.700 1359.140 2934.200 1362.140 ;
        RECT -14.580 1359.130 -11.580 1359.140 ;
        RECT 2931.200 1359.130 2934.200 1359.140 ;
        RECT -14.580 1182.140 -11.580 1182.150 ;
        RECT 2931.200 1182.140 2934.200 1182.150 ;
        RECT -14.580 1179.140 0.300 1182.140 ;
        RECT 2919.700 1179.140 2934.200 1182.140 ;
        RECT -14.580 1179.130 -11.580 1179.140 ;
        RECT 2931.200 1179.130 2934.200 1179.140 ;
        RECT -14.580 1002.140 -11.580 1002.150 ;
        RECT 2931.200 1002.140 2934.200 1002.150 ;
        RECT -14.580 999.140 0.300 1002.140 ;
        RECT 2919.700 999.140 2934.200 1002.140 ;
        RECT -14.580 999.130 -11.580 999.140 ;
        RECT 2931.200 999.130 2934.200 999.140 ;
        RECT -14.580 822.140 -11.580 822.150 ;
        RECT 2931.200 822.140 2934.200 822.150 ;
        RECT -14.580 819.140 0.300 822.140 ;
        RECT 2919.700 819.140 2934.200 822.140 ;
        RECT -14.580 819.130 -11.580 819.140 ;
        RECT 2931.200 819.130 2934.200 819.140 ;
        RECT -14.580 642.140 -11.580 642.150 ;
        RECT 2931.200 642.140 2934.200 642.150 ;
        RECT -14.580 639.140 0.300 642.140 ;
        RECT 2919.700 639.140 2934.200 642.140 ;
        RECT -14.580 639.130 -11.580 639.140 ;
        RECT 2931.200 639.130 2934.200 639.140 ;
        RECT -14.580 462.140 -11.580 462.150 ;
        RECT 2931.200 462.140 2934.200 462.150 ;
        RECT -14.580 459.140 0.300 462.140 ;
        RECT 2919.700 459.140 2934.200 462.140 ;
        RECT -14.580 459.130 -11.580 459.140 ;
        RECT 2931.200 459.130 2934.200 459.140 ;
        RECT -14.580 282.140 -11.580 282.150 ;
        RECT 2931.200 282.140 2934.200 282.150 ;
        RECT -14.580 279.140 0.300 282.140 ;
        RECT 2919.700 279.140 2934.200 282.140 ;
        RECT -14.580 279.130 -11.580 279.140 ;
        RECT 2931.200 279.130 2934.200 279.140 ;
        RECT -14.580 102.140 -11.580 102.150 ;
        RECT 2931.200 102.140 2934.200 102.150 ;
        RECT -14.580 99.140 0.300 102.140 ;
        RECT 2919.700 99.140 2934.200 102.140 ;
        RECT -14.580 99.130 -11.580 99.140 ;
        RECT 2931.200 99.130 2934.200 99.140 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 3519.700 25.020 3538.100 ;
        RECT 202.020 3519.700 205.020 3538.100 ;
        RECT 382.020 3519.700 385.020 3538.100 ;
        RECT 562.020 3519.700 565.020 3538.100 ;
        RECT 742.020 3519.700 745.020 3538.100 ;
        RECT 922.020 3519.700 925.020 3538.100 ;
        RECT 1102.020 3519.700 1105.020 3538.100 ;
        RECT 1282.020 3519.700 1285.020 3538.100 ;
        RECT 1462.020 3519.700 1465.020 3538.100 ;
        RECT 1642.020 3519.700 1645.020 3538.100 ;
        RECT 1822.020 3519.700 1825.020 3538.100 ;
        RECT 2002.020 3519.700 2005.020 3538.100 ;
        RECT 2182.020 3519.700 2185.020 3538.100 ;
        RECT 2362.020 3519.700 2365.020 3538.100 ;
        RECT 2542.020 3519.700 2545.020 3538.100 ;
        RECT 2722.020 3519.700 2725.020 3538.100 ;
        RECT 2902.020 3519.700 2905.020 3538.100 ;
        RECT 22.020 -18.420 25.020 0.300 ;
        RECT 202.020 -18.420 205.020 0.300 ;
        RECT 382.020 -18.420 385.020 0.300 ;
        RECT 562.020 -18.420 565.020 0.300 ;
        RECT 742.020 -18.420 745.020 0.300 ;
        RECT 922.020 -18.420 925.020 0.300 ;
        RECT 1102.020 -18.420 1105.020 0.300 ;
        RECT 1282.020 -18.420 1285.020 0.300 ;
        RECT 1462.020 -18.420 1465.020 0.300 ;
        RECT 1642.020 -18.420 1645.020 0.300 ;
        RECT 1822.020 -18.420 1825.020 0.300 ;
        RECT 2002.020 -18.420 2005.020 0.300 ;
        RECT 2182.020 -18.420 2185.020 0.300 ;
        RECT 2362.020 -18.420 2365.020 0.300 ;
        RECT 2542.020 -18.420 2545.020 0.300 ;
        RECT 2722.020 -18.420 2725.020 0.300 ;
        RECT 2902.020 -18.420 2905.020 0.300 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT -18.270 3448.850 -17.090 3450.030 ;
        RECT -18.270 3447.250 -17.090 3448.430 ;
        RECT -18.270 3268.850 -17.090 3270.030 ;
        RECT -18.270 3267.250 -17.090 3268.430 ;
        RECT -18.270 3088.850 -17.090 3090.030 ;
        RECT -18.270 3087.250 -17.090 3088.430 ;
        RECT -18.270 2908.850 -17.090 2910.030 ;
        RECT -18.270 2907.250 -17.090 2908.430 ;
        RECT -18.270 2728.850 -17.090 2730.030 ;
        RECT -18.270 2727.250 -17.090 2728.430 ;
        RECT -18.270 2548.850 -17.090 2550.030 ;
        RECT -18.270 2547.250 -17.090 2548.430 ;
        RECT -18.270 2368.850 -17.090 2370.030 ;
        RECT -18.270 2367.250 -17.090 2368.430 ;
        RECT -18.270 2188.850 -17.090 2190.030 ;
        RECT -18.270 2187.250 -17.090 2188.430 ;
        RECT -18.270 2008.850 -17.090 2010.030 ;
        RECT -18.270 2007.250 -17.090 2008.430 ;
        RECT -18.270 1828.850 -17.090 1830.030 ;
        RECT -18.270 1827.250 -17.090 1828.430 ;
        RECT -18.270 1648.850 -17.090 1650.030 ;
        RECT -18.270 1647.250 -17.090 1648.430 ;
        RECT -18.270 1468.850 -17.090 1470.030 ;
        RECT -18.270 1467.250 -17.090 1468.430 ;
        RECT -18.270 1288.850 -17.090 1290.030 ;
        RECT -18.270 1287.250 -17.090 1288.430 ;
        RECT -18.270 1108.850 -17.090 1110.030 ;
        RECT -18.270 1107.250 -17.090 1108.430 ;
        RECT -18.270 928.850 -17.090 930.030 ;
        RECT -18.270 927.250 -17.090 928.430 ;
        RECT -18.270 748.850 -17.090 750.030 ;
        RECT -18.270 747.250 -17.090 748.430 ;
        RECT -18.270 568.850 -17.090 570.030 ;
        RECT -18.270 567.250 -17.090 568.430 ;
        RECT -18.270 388.850 -17.090 390.030 ;
        RECT -18.270 387.250 -17.090 388.430 ;
        RECT -18.270 208.850 -17.090 210.030 ;
        RECT -18.270 207.250 -17.090 208.430 ;
        RECT -18.270 28.850 -17.090 30.030 ;
        RECT -18.270 27.250 -17.090 28.430 ;
        RECT 2936.710 3448.850 2937.890 3450.030 ;
        RECT 2936.710 3447.250 2937.890 3448.430 ;
        RECT 2936.710 3268.850 2937.890 3270.030 ;
        RECT 2936.710 3267.250 2937.890 3268.430 ;
        RECT 2936.710 3088.850 2937.890 3090.030 ;
        RECT 2936.710 3087.250 2937.890 3088.430 ;
        RECT 2936.710 2908.850 2937.890 2910.030 ;
        RECT 2936.710 2907.250 2937.890 2908.430 ;
        RECT 2936.710 2728.850 2937.890 2730.030 ;
        RECT 2936.710 2727.250 2937.890 2728.430 ;
        RECT 2936.710 2548.850 2937.890 2550.030 ;
        RECT 2936.710 2547.250 2937.890 2548.430 ;
        RECT 2936.710 2368.850 2937.890 2370.030 ;
        RECT 2936.710 2367.250 2937.890 2368.430 ;
        RECT 2936.710 2188.850 2937.890 2190.030 ;
        RECT 2936.710 2187.250 2937.890 2188.430 ;
        RECT 2936.710 2008.850 2937.890 2010.030 ;
        RECT 2936.710 2007.250 2937.890 2008.430 ;
        RECT 2936.710 1828.850 2937.890 1830.030 ;
        RECT 2936.710 1827.250 2937.890 1828.430 ;
        RECT 2936.710 1648.850 2937.890 1650.030 ;
        RECT 2936.710 1647.250 2937.890 1648.430 ;
        RECT 2936.710 1468.850 2937.890 1470.030 ;
        RECT 2936.710 1467.250 2937.890 1468.430 ;
        RECT 2936.710 1288.850 2937.890 1290.030 ;
        RECT 2936.710 1287.250 2937.890 1288.430 ;
        RECT 2936.710 1108.850 2937.890 1110.030 ;
        RECT 2936.710 1107.250 2937.890 1108.430 ;
        RECT 2936.710 928.850 2937.890 930.030 ;
        RECT 2936.710 927.250 2937.890 928.430 ;
        RECT 2936.710 748.850 2937.890 750.030 ;
        RECT 2936.710 747.250 2937.890 748.430 ;
        RECT 2936.710 568.850 2937.890 570.030 ;
        RECT 2936.710 567.250 2937.890 568.430 ;
        RECT 2936.710 388.850 2937.890 390.030 ;
        RECT 2936.710 387.250 2937.890 388.430 ;
        RECT 2936.710 208.850 2937.890 210.030 ;
        RECT 2936.710 207.250 2937.890 208.430 ;
        RECT 2936.710 28.850 2937.890 30.030 ;
        RECT 2936.710 27.250 2937.890 28.430 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.140 -16.180 3450.150 ;
        RECT 2935.800 3450.140 2938.800 3450.150 ;
        RECT -23.780 3447.140 0.300 3450.140 ;
        RECT 2919.700 3447.140 2943.400 3450.140 ;
        RECT -19.180 3447.130 -16.180 3447.140 ;
        RECT 2935.800 3447.130 2938.800 3447.140 ;
        RECT -19.180 3270.140 -16.180 3270.150 ;
        RECT 2935.800 3270.140 2938.800 3270.150 ;
        RECT -23.780 3267.140 0.300 3270.140 ;
        RECT 2919.700 3267.140 2943.400 3270.140 ;
        RECT -19.180 3267.130 -16.180 3267.140 ;
        RECT 2935.800 3267.130 2938.800 3267.140 ;
        RECT -19.180 3090.140 -16.180 3090.150 ;
        RECT 2935.800 3090.140 2938.800 3090.150 ;
        RECT -23.780 3087.140 0.300 3090.140 ;
        RECT 2919.700 3087.140 2943.400 3090.140 ;
        RECT -19.180 3087.130 -16.180 3087.140 ;
        RECT 2935.800 3087.130 2938.800 3087.140 ;
        RECT -19.180 2910.140 -16.180 2910.150 ;
        RECT 2935.800 2910.140 2938.800 2910.150 ;
        RECT -23.780 2907.140 0.300 2910.140 ;
        RECT 2919.700 2907.140 2943.400 2910.140 ;
        RECT -19.180 2907.130 -16.180 2907.140 ;
        RECT 2935.800 2907.130 2938.800 2907.140 ;
        RECT -19.180 2730.140 -16.180 2730.150 ;
        RECT 2935.800 2730.140 2938.800 2730.150 ;
        RECT -23.780 2727.140 0.300 2730.140 ;
        RECT 2919.700 2727.140 2943.400 2730.140 ;
        RECT -19.180 2727.130 -16.180 2727.140 ;
        RECT 2935.800 2727.130 2938.800 2727.140 ;
        RECT -19.180 2550.140 -16.180 2550.150 ;
        RECT 2935.800 2550.140 2938.800 2550.150 ;
        RECT -23.780 2547.140 0.300 2550.140 ;
        RECT 2919.700 2547.140 2943.400 2550.140 ;
        RECT -19.180 2547.130 -16.180 2547.140 ;
        RECT 2935.800 2547.130 2938.800 2547.140 ;
        RECT -19.180 2370.140 -16.180 2370.150 ;
        RECT 2935.800 2370.140 2938.800 2370.150 ;
        RECT -23.780 2367.140 0.300 2370.140 ;
        RECT 2919.700 2367.140 2943.400 2370.140 ;
        RECT -19.180 2367.130 -16.180 2367.140 ;
        RECT 2935.800 2367.130 2938.800 2367.140 ;
        RECT -19.180 2190.140 -16.180 2190.150 ;
        RECT 2935.800 2190.140 2938.800 2190.150 ;
        RECT -23.780 2187.140 0.300 2190.140 ;
        RECT 2919.700 2187.140 2943.400 2190.140 ;
        RECT -19.180 2187.130 -16.180 2187.140 ;
        RECT 2935.800 2187.130 2938.800 2187.140 ;
        RECT -19.180 2010.140 -16.180 2010.150 ;
        RECT 2935.800 2010.140 2938.800 2010.150 ;
        RECT -23.780 2007.140 0.300 2010.140 ;
        RECT 2919.700 2007.140 2943.400 2010.140 ;
        RECT -19.180 2007.130 -16.180 2007.140 ;
        RECT 2935.800 2007.130 2938.800 2007.140 ;
        RECT -19.180 1830.140 -16.180 1830.150 ;
        RECT 2935.800 1830.140 2938.800 1830.150 ;
        RECT -23.780 1827.140 0.300 1830.140 ;
        RECT 2919.700 1827.140 2943.400 1830.140 ;
        RECT -19.180 1827.130 -16.180 1827.140 ;
        RECT 2935.800 1827.130 2938.800 1827.140 ;
        RECT -19.180 1650.140 -16.180 1650.150 ;
        RECT 2935.800 1650.140 2938.800 1650.150 ;
        RECT -23.780 1647.140 0.300 1650.140 ;
        RECT 2919.700 1647.140 2943.400 1650.140 ;
        RECT -19.180 1647.130 -16.180 1647.140 ;
        RECT 2935.800 1647.130 2938.800 1647.140 ;
        RECT -19.180 1470.140 -16.180 1470.150 ;
        RECT 2935.800 1470.140 2938.800 1470.150 ;
        RECT -23.780 1467.140 0.300 1470.140 ;
        RECT 2919.700 1467.140 2943.400 1470.140 ;
        RECT -19.180 1467.130 -16.180 1467.140 ;
        RECT 2935.800 1467.130 2938.800 1467.140 ;
        RECT -19.180 1290.140 -16.180 1290.150 ;
        RECT 2935.800 1290.140 2938.800 1290.150 ;
        RECT -23.780 1287.140 0.300 1290.140 ;
        RECT 2919.700 1287.140 2943.400 1290.140 ;
        RECT -19.180 1287.130 -16.180 1287.140 ;
        RECT 2935.800 1287.130 2938.800 1287.140 ;
        RECT -19.180 1110.140 -16.180 1110.150 ;
        RECT 2935.800 1110.140 2938.800 1110.150 ;
        RECT -23.780 1107.140 0.300 1110.140 ;
        RECT 2919.700 1107.140 2943.400 1110.140 ;
        RECT -19.180 1107.130 -16.180 1107.140 ;
        RECT 2935.800 1107.130 2938.800 1107.140 ;
        RECT -19.180 930.140 -16.180 930.150 ;
        RECT 2935.800 930.140 2938.800 930.150 ;
        RECT -23.780 927.140 0.300 930.140 ;
        RECT 2919.700 927.140 2943.400 930.140 ;
        RECT -19.180 927.130 -16.180 927.140 ;
        RECT 2935.800 927.130 2938.800 927.140 ;
        RECT -19.180 750.140 -16.180 750.150 ;
        RECT 2935.800 750.140 2938.800 750.150 ;
        RECT -23.780 747.140 0.300 750.140 ;
        RECT 2919.700 747.140 2943.400 750.140 ;
        RECT -19.180 747.130 -16.180 747.140 ;
        RECT 2935.800 747.130 2938.800 747.140 ;
        RECT -19.180 570.140 -16.180 570.150 ;
        RECT 2935.800 570.140 2938.800 570.150 ;
        RECT -23.780 567.140 0.300 570.140 ;
        RECT 2919.700 567.140 2943.400 570.140 ;
        RECT -19.180 567.130 -16.180 567.140 ;
        RECT 2935.800 567.130 2938.800 567.140 ;
        RECT -19.180 390.140 -16.180 390.150 ;
        RECT 2935.800 390.140 2938.800 390.150 ;
        RECT -23.780 387.140 0.300 390.140 ;
        RECT 2919.700 387.140 2943.400 390.140 ;
        RECT -19.180 387.130 -16.180 387.140 ;
        RECT 2935.800 387.130 2938.800 387.140 ;
        RECT -19.180 210.140 -16.180 210.150 ;
        RECT 2935.800 210.140 2938.800 210.150 ;
        RECT -23.780 207.140 0.300 210.140 ;
        RECT 2919.700 207.140 2943.400 210.140 ;
        RECT -19.180 207.130 -16.180 207.140 ;
        RECT 2935.800 207.130 2938.800 207.140 ;
        RECT -19.180 30.140 -16.180 30.150 ;
        RECT 2935.800 30.140 2938.800 30.150 ;
        RECT -23.780 27.140 0.300 30.140 ;
        RECT 2919.700 27.140 2943.400 30.140 ;
        RECT -19.180 27.130 -16.180 27.140 ;
        RECT 2935.800 27.130 2938.800 27.140 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 3519.700 115.020 3538.100 ;
        RECT 292.020 3519.700 295.020 3538.100 ;
        RECT 472.020 3519.700 475.020 3538.100 ;
        RECT 652.020 3519.700 655.020 3538.100 ;
        RECT 832.020 3519.700 835.020 3538.100 ;
        RECT 1012.020 3519.700 1015.020 3538.100 ;
        RECT 1192.020 3519.700 1195.020 3538.100 ;
        RECT 1372.020 3519.700 1375.020 3538.100 ;
        RECT 1552.020 3519.700 1555.020 3538.100 ;
        RECT 1732.020 3519.700 1735.020 3538.100 ;
        RECT 1912.020 3519.700 1915.020 3538.100 ;
        RECT 2092.020 3519.700 2095.020 3538.100 ;
        RECT 2272.020 3519.700 2275.020 3538.100 ;
        RECT 2452.020 3519.700 2455.020 3538.100 ;
        RECT 2632.020 3519.700 2635.020 3538.100 ;
        RECT 2812.020 3519.700 2815.020 3538.100 ;
        RECT 112.020 -18.420 115.020 0.300 ;
        RECT 292.020 -18.420 295.020 0.300 ;
        RECT 472.020 -18.420 475.020 0.300 ;
        RECT 652.020 -18.420 655.020 0.300 ;
        RECT 832.020 -18.420 835.020 0.300 ;
        RECT 1012.020 -18.420 1015.020 0.300 ;
        RECT 1192.020 -18.420 1195.020 0.300 ;
        RECT 1372.020 -18.420 1375.020 0.300 ;
        RECT 1552.020 -18.420 1555.020 0.300 ;
        RECT 1732.020 -18.420 1735.020 0.300 ;
        RECT 1912.020 -18.420 1915.020 0.300 ;
        RECT 2092.020 -18.420 2095.020 0.300 ;
        RECT 2272.020 -18.420 2275.020 0.300 ;
        RECT 2452.020 -18.420 2455.020 0.300 ;
        RECT 2632.020 -18.420 2635.020 0.300 ;
        RECT 2812.020 -18.420 2815.020 0.300 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT -22.870 3358.850 -21.690 3360.030 ;
        RECT -22.870 3357.250 -21.690 3358.430 ;
        RECT -22.870 3178.850 -21.690 3180.030 ;
        RECT -22.870 3177.250 -21.690 3178.430 ;
        RECT -22.870 2998.850 -21.690 3000.030 ;
        RECT -22.870 2997.250 -21.690 2998.430 ;
        RECT -22.870 2818.850 -21.690 2820.030 ;
        RECT -22.870 2817.250 -21.690 2818.430 ;
        RECT -22.870 2638.850 -21.690 2640.030 ;
        RECT -22.870 2637.250 -21.690 2638.430 ;
        RECT -22.870 2458.850 -21.690 2460.030 ;
        RECT -22.870 2457.250 -21.690 2458.430 ;
        RECT -22.870 2278.850 -21.690 2280.030 ;
        RECT -22.870 2277.250 -21.690 2278.430 ;
        RECT -22.870 2098.850 -21.690 2100.030 ;
        RECT -22.870 2097.250 -21.690 2098.430 ;
        RECT -22.870 1918.850 -21.690 1920.030 ;
        RECT -22.870 1917.250 -21.690 1918.430 ;
        RECT -22.870 1738.850 -21.690 1740.030 ;
        RECT -22.870 1737.250 -21.690 1738.430 ;
        RECT -22.870 1558.850 -21.690 1560.030 ;
        RECT -22.870 1557.250 -21.690 1558.430 ;
        RECT -22.870 1378.850 -21.690 1380.030 ;
        RECT -22.870 1377.250 -21.690 1378.430 ;
        RECT -22.870 1198.850 -21.690 1200.030 ;
        RECT -22.870 1197.250 -21.690 1198.430 ;
        RECT -22.870 1018.850 -21.690 1020.030 ;
        RECT -22.870 1017.250 -21.690 1018.430 ;
        RECT -22.870 838.850 -21.690 840.030 ;
        RECT -22.870 837.250 -21.690 838.430 ;
        RECT -22.870 658.850 -21.690 660.030 ;
        RECT -22.870 657.250 -21.690 658.430 ;
        RECT -22.870 478.850 -21.690 480.030 ;
        RECT -22.870 477.250 -21.690 478.430 ;
        RECT -22.870 298.850 -21.690 300.030 ;
        RECT -22.870 297.250 -21.690 298.430 ;
        RECT -22.870 118.850 -21.690 120.030 ;
        RECT -22.870 117.250 -21.690 118.430 ;
        RECT 2941.310 3358.850 2942.490 3360.030 ;
        RECT 2941.310 3357.250 2942.490 3358.430 ;
        RECT 2941.310 3178.850 2942.490 3180.030 ;
        RECT 2941.310 3177.250 2942.490 3178.430 ;
        RECT 2941.310 2998.850 2942.490 3000.030 ;
        RECT 2941.310 2997.250 2942.490 2998.430 ;
        RECT 2941.310 2818.850 2942.490 2820.030 ;
        RECT 2941.310 2817.250 2942.490 2818.430 ;
        RECT 2941.310 2638.850 2942.490 2640.030 ;
        RECT 2941.310 2637.250 2942.490 2638.430 ;
        RECT 2941.310 2458.850 2942.490 2460.030 ;
        RECT 2941.310 2457.250 2942.490 2458.430 ;
        RECT 2941.310 2278.850 2942.490 2280.030 ;
        RECT 2941.310 2277.250 2942.490 2278.430 ;
        RECT 2941.310 2098.850 2942.490 2100.030 ;
        RECT 2941.310 2097.250 2942.490 2098.430 ;
        RECT 2941.310 1918.850 2942.490 1920.030 ;
        RECT 2941.310 1917.250 2942.490 1918.430 ;
        RECT 2941.310 1738.850 2942.490 1740.030 ;
        RECT 2941.310 1737.250 2942.490 1738.430 ;
        RECT 2941.310 1558.850 2942.490 1560.030 ;
        RECT 2941.310 1557.250 2942.490 1558.430 ;
        RECT 2941.310 1378.850 2942.490 1380.030 ;
        RECT 2941.310 1377.250 2942.490 1378.430 ;
        RECT 2941.310 1198.850 2942.490 1200.030 ;
        RECT 2941.310 1197.250 2942.490 1198.430 ;
        RECT 2941.310 1018.850 2942.490 1020.030 ;
        RECT 2941.310 1017.250 2942.490 1018.430 ;
        RECT 2941.310 838.850 2942.490 840.030 ;
        RECT 2941.310 837.250 2942.490 838.430 ;
        RECT 2941.310 658.850 2942.490 660.030 ;
        RECT 2941.310 657.250 2942.490 658.430 ;
        RECT 2941.310 478.850 2942.490 480.030 ;
        RECT 2941.310 477.250 2942.490 478.430 ;
        RECT 2941.310 298.850 2942.490 300.030 ;
        RECT 2941.310 297.250 2942.490 298.430 ;
        RECT 2941.310 118.850 2942.490 120.030 ;
        RECT 2941.310 117.250 2942.490 118.430 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.140 -20.780 3360.150 ;
        RECT 2940.400 3360.140 2943.400 3360.150 ;
        RECT -23.780 3357.140 0.300 3360.140 ;
        RECT 2919.700 3357.140 2943.400 3360.140 ;
        RECT -23.780 3357.130 -20.780 3357.140 ;
        RECT 2940.400 3357.130 2943.400 3357.140 ;
        RECT -23.780 3180.140 -20.780 3180.150 ;
        RECT 2940.400 3180.140 2943.400 3180.150 ;
        RECT -23.780 3177.140 0.300 3180.140 ;
        RECT 2919.700 3177.140 2943.400 3180.140 ;
        RECT -23.780 3177.130 -20.780 3177.140 ;
        RECT 2940.400 3177.130 2943.400 3177.140 ;
        RECT -23.780 3000.140 -20.780 3000.150 ;
        RECT 2940.400 3000.140 2943.400 3000.150 ;
        RECT -23.780 2997.140 0.300 3000.140 ;
        RECT 2919.700 2997.140 2943.400 3000.140 ;
        RECT -23.780 2997.130 -20.780 2997.140 ;
        RECT 2940.400 2997.130 2943.400 2997.140 ;
        RECT -23.780 2820.140 -20.780 2820.150 ;
        RECT 2940.400 2820.140 2943.400 2820.150 ;
        RECT -23.780 2817.140 0.300 2820.140 ;
        RECT 2919.700 2817.140 2943.400 2820.140 ;
        RECT -23.780 2817.130 -20.780 2817.140 ;
        RECT 2940.400 2817.130 2943.400 2817.140 ;
        RECT -23.780 2640.140 -20.780 2640.150 ;
        RECT 2940.400 2640.140 2943.400 2640.150 ;
        RECT -23.780 2637.140 0.300 2640.140 ;
        RECT 2919.700 2637.140 2943.400 2640.140 ;
        RECT -23.780 2637.130 -20.780 2637.140 ;
        RECT 2940.400 2637.130 2943.400 2637.140 ;
        RECT -23.780 2460.140 -20.780 2460.150 ;
        RECT 2940.400 2460.140 2943.400 2460.150 ;
        RECT -23.780 2457.140 0.300 2460.140 ;
        RECT 2919.700 2457.140 2943.400 2460.140 ;
        RECT -23.780 2457.130 -20.780 2457.140 ;
        RECT 2940.400 2457.130 2943.400 2457.140 ;
        RECT -23.780 2280.140 -20.780 2280.150 ;
        RECT 2940.400 2280.140 2943.400 2280.150 ;
        RECT -23.780 2277.140 0.300 2280.140 ;
        RECT 2919.700 2277.140 2943.400 2280.140 ;
        RECT -23.780 2277.130 -20.780 2277.140 ;
        RECT 2940.400 2277.130 2943.400 2277.140 ;
        RECT -23.780 2100.140 -20.780 2100.150 ;
        RECT 2940.400 2100.140 2943.400 2100.150 ;
        RECT -23.780 2097.140 0.300 2100.140 ;
        RECT 2919.700 2097.140 2943.400 2100.140 ;
        RECT -23.780 2097.130 -20.780 2097.140 ;
        RECT 2940.400 2097.130 2943.400 2097.140 ;
        RECT -23.780 1920.140 -20.780 1920.150 ;
        RECT 2940.400 1920.140 2943.400 1920.150 ;
        RECT -23.780 1917.140 0.300 1920.140 ;
        RECT 2919.700 1917.140 2943.400 1920.140 ;
        RECT -23.780 1917.130 -20.780 1917.140 ;
        RECT 2940.400 1917.130 2943.400 1917.140 ;
        RECT -23.780 1740.140 -20.780 1740.150 ;
        RECT 2940.400 1740.140 2943.400 1740.150 ;
        RECT -23.780 1737.140 0.300 1740.140 ;
        RECT 2919.700 1737.140 2943.400 1740.140 ;
        RECT -23.780 1737.130 -20.780 1737.140 ;
        RECT 2940.400 1737.130 2943.400 1737.140 ;
        RECT -23.780 1560.140 -20.780 1560.150 ;
        RECT 2940.400 1560.140 2943.400 1560.150 ;
        RECT -23.780 1557.140 0.300 1560.140 ;
        RECT 2919.700 1557.140 2943.400 1560.140 ;
        RECT -23.780 1557.130 -20.780 1557.140 ;
        RECT 2940.400 1557.130 2943.400 1557.140 ;
        RECT -23.780 1380.140 -20.780 1380.150 ;
        RECT 2940.400 1380.140 2943.400 1380.150 ;
        RECT -23.780 1377.140 0.300 1380.140 ;
        RECT 2919.700 1377.140 2943.400 1380.140 ;
        RECT -23.780 1377.130 -20.780 1377.140 ;
        RECT 2940.400 1377.130 2943.400 1377.140 ;
        RECT -23.780 1200.140 -20.780 1200.150 ;
        RECT 2940.400 1200.140 2943.400 1200.150 ;
        RECT -23.780 1197.140 0.300 1200.140 ;
        RECT 2919.700 1197.140 2943.400 1200.140 ;
        RECT -23.780 1197.130 -20.780 1197.140 ;
        RECT 2940.400 1197.130 2943.400 1197.140 ;
        RECT -23.780 1020.140 -20.780 1020.150 ;
        RECT 2940.400 1020.140 2943.400 1020.150 ;
        RECT -23.780 1017.140 0.300 1020.140 ;
        RECT 2919.700 1017.140 2943.400 1020.140 ;
        RECT -23.780 1017.130 -20.780 1017.140 ;
        RECT 2940.400 1017.130 2943.400 1017.140 ;
        RECT -23.780 840.140 -20.780 840.150 ;
        RECT 2940.400 840.140 2943.400 840.150 ;
        RECT -23.780 837.140 0.300 840.140 ;
        RECT 2919.700 837.140 2943.400 840.140 ;
        RECT -23.780 837.130 -20.780 837.140 ;
        RECT 2940.400 837.130 2943.400 837.140 ;
        RECT -23.780 660.140 -20.780 660.150 ;
        RECT 2940.400 660.140 2943.400 660.150 ;
        RECT -23.780 657.140 0.300 660.140 ;
        RECT 2919.700 657.140 2943.400 660.140 ;
        RECT -23.780 657.130 -20.780 657.140 ;
        RECT 2940.400 657.130 2943.400 657.140 ;
        RECT -23.780 480.140 -20.780 480.150 ;
        RECT 2940.400 480.140 2943.400 480.150 ;
        RECT -23.780 477.140 0.300 480.140 ;
        RECT 2919.700 477.140 2943.400 480.140 ;
        RECT -23.780 477.130 -20.780 477.140 ;
        RECT 2940.400 477.130 2943.400 477.140 ;
        RECT -23.780 300.140 -20.780 300.150 ;
        RECT 2940.400 300.140 2943.400 300.150 ;
        RECT -23.780 297.140 0.300 300.140 ;
        RECT 2919.700 297.140 2943.400 300.140 ;
        RECT -23.780 297.130 -20.780 297.140 ;
        RECT 2940.400 297.130 2943.400 297.140 ;
        RECT -23.780 120.140 -20.780 120.150 ;
        RECT 2940.400 120.140 2943.400 120.150 ;
        RECT -23.780 117.140 0.300 120.140 ;
        RECT 2919.700 117.140 2943.400 120.140 ;
        RECT -23.780 117.130 -20.780 117.140 ;
        RECT 2940.400 117.130 2943.400 117.140 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 3519.700 43.020 3547.300 ;
        RECT 220.020 3519.700 223.020 3547.300 ;
        RECT 400.020 3519.700 403.020 3547.300 ;
        RECT 580.020 3519.700 583.020 3547.300 ;
        RECT 760.020 3519.700 763.020 3547.300 ;
        RECT 940.020 3519.700 943.020 3547.300 ;
        RECT 1120.020 3519.700 1123.020 3547.300 ;
        RECT 1300.020 3519.700 1303.020 3547.300 ;
        RECT 1480.020 3519.700 1483.020 3547.300 ;
        RECT 1660.020 3519.700 1663.020 3547.300 ;
        RECT 1840.020 3519.700 1843.020 3547.300 ;
        RECT 2020.020 3519.700 2023.020 3547.300 ;
        RECT 2200.020 3519.700 2203.020 3547.300 ;
        RECT 2380.020 3519.700 2383.020 3547.300 ;
        RECT 2560.020 3519.700 2563.020 3547.300 ;
        RECT 2740.020 3519.700 2743.020 3547.300 ;
        RECT 40.020 -27.620 43.020 0.300 ;
        RECT 220.020 -27.620 223.020 0.300 ;
        RECT 400.020 -27.620 403.020 0.300 ;
        RECT 580.020 -27.620 583.020 0.300 ;
        RECT 760.020 -27.620 763.020 0.300 ;
        RECT 940.020 -27.620 943.020 0.300 ;
        RECT 1120.020 -27.620 1123.020 0.300 ;
        RECT 1300.020 -27.620 1303.020 0.300 ;
        RECT 1480.020 -27.620 1483.020 0.300 ;
        RECT 1660.020 -27.620 1663.020 0.300 ;
        RECT 1840.020 -27.620 1843.020 0.300 ;
        RECT 2020.020 -27.620 2023.020 0.300 ;
        RECT 2200.020 -27.620 2203.020 0.300 ;
        RECT 2380.020 -27.620 2383.020 0.300 ;
        RECT 2560.020 -27.620 2563.020 0.300 ;
        RECT 2740.020 -27.620 2743.020 0.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT -27.470 3466.850 -26.290 3468.030 ;
        RECT -27.470 3465.250 -26.290 3466.430 ;
        RECT -27.470 3286.850 -26.290 3288.030 ;
        RECT -27.470 3285.250 -26.290 3286.430 ;
        RECT -27.470 3106.850 -26.290 3108.030 ;
        RECT -27.470 3105.250 -26.290 3106.430 ;
        RECT -27.470 2926.850 -26.290 2928.030 ;
        RECT -27.470 2925.250 -26.290 2926.430 ;
        RECT -27.470 2746.850 -26.290 2748.030 ;
        RECT -27.470 2745.250 -26.290 2746.430 ;
        RECT -27.470 2566.850 -26.290 2568.030 ;
        RECT -27.470 2565.250 -26.290 2566.430 ;
        RECT -27.470 2386.850 -26.290 2388.030 ;
        RECT -27.470 2385.250 -26.290 2386.430 ;
        RECT -27.470 2206.850 -26.290 2208.030 ;
        RECT -27.470 2205.250 -26.290 2206.430 ;
        RECT -27.470 2026.850 -26.290 2028.030 ;
        RECT -27.470 2025.250 -26.290 2026.430 ;
        RECT -27.470 1846.850 -26.290 1848.030 ;
        RECT -27.470 1845.250 -26.290 1846.430 ;
        RECT -27.470 1666.850 -26.290 1668.030 ;
        RECT -27.470 1665.250 -26.290 1666.430 ;
        RECT -27.470 1486.850 -26.290 1488.030 ;
        RECT -27.470 1485.250 -26.290 1486.430 ;
        RECT -27.470 1306.850 -26.290 1308.030 ;
        RECT -27.470 1305.250 -26.290 1306.430 ;
        RECT -27.470 1126.850 -26.290 1128.030 ;
        RECT -27.470 1125.250 -26.290 1126.430 ;
        RECT -27.470 946.850 -26.290 948.030 ;
        RECT -27.470 945.250 -26.290 946.430 ;
        RECT -27.470 766.850 -26.290 768.030 ;
        RECT -27.470 765.250 -26.290 766.430 ;
        RECT -27.470 586.850 -26.290 588.030 ;
        RECT -27.470 585.250 -26.290 586.430 ;
        RECT -27.470 406.850 -26.290 408.030 ;
        RECT -27.470 405.250 -26.290 406.430 ;
        RECT -27.470 226.850 -26.290 228.030 ;
        RECT -27.470 225.250 -26.290 226.430 ;
        RECT -27.470 46.850 -26.290 48.030 ;
        RECT -27.470 45.250 -26.290 46.430 ;
        RECT 2945.910 3466.850 2947.090 3468.030 ;
        RECT 2945.910 3465.250 2947.090 3466.430 ;
        RECT 2945.910 3286.850 2947.090 3288.030 ;
        RECT 2945.910 3285.250 2947.090 3286.430 ;
        RECT 2945.910 3106.850 2947.090 3108.030 ;
        RECT 2945.910 3105.250 2947.090 3106.430 ;
        RECT 2945.910 2926.850 2947.090 2928.030 ;
        RECT 2945.910 2925.250 2947.090 2926.430 ;
        RECT 2945.910 2746.850 2947.090 2748.030 ;
        RECT 2945.910 2745.250 2947.090 2746.430 ;
        RECT 2945.910 2566.850 2947.090 2568.030 ;
        RECT 2945.910 2565.250 2947.090 2566.430 ;
        RECT 2945.910 2386.850 2947.090 2388.030 ;
        RECT 2945.910 2385.250 2947.090 2386.430 ;
        RECT 2945.910 2206.850 2947.090 2208.030 ;
        RECT 2945.910 2205.250 2947.090 2206.430 ;
        RECT 2945.910 2026.850 2947.090 2028.030 ;
        RECT 2945.910 2025.250 2947.090 2026.430 ;
        RECT 2945.910 1846.850 2947.090 1848.030 ;
        RECT 2945.910 1845.250 2947.090 1846.430 ;
        RECT 2945.910 1666.850 2947.090 1668.030 ;
        RECT 2945.910 1665.250 2947.090 1666.430 ;
        RECT 2945.910 1486.850 2947.090 1488.030 ;
        RECT 2945.910 1485.250 2947.090 1486.430 ;
        RECT 2945.910 1306.850 2947.090 1308.030 ;
        RECT 2945.910 1305.250 2947.090 1306.430 ;
        RECT 2945.910 1126.850 2947.090 1128.030 ;
        RECT 2945.910 1125.250 2947.090 1126.430 ;
        RECT 2945.910 946.850 2947.090 948.030 ;
        RECT 2945.910 945.250 2947.090 946.430 ;
        RECT 2945.910 766.850 2947.090 768.030 ;
        RECT 2945.910 765.250 2947.090 766.430 ;
        RECT 2945.910 586.850 2947.090 588.030 ;
        RECT 2945.910 585.250 2947.090 586.430 ;
        RECT 2945.910 406.850 2947.090 408.030 ;
        RECT 2945.910 405.250 2947.090 406.430 ;
        RECT 2945.910 226.850 2947.090 228.030 ;
        RECT 2945.910 225.250 2947.090 226.430 ;
        RECT 2945.910 46.850 2947.090 48.030 ;
        RECT 2945.910 45.250 2947.090 46.430 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.140 -25.380 3468.150 ;
        RECT 2945.000 3468.140 2948.000 3468.150 ;
        RECT -32.980 3465.140 0.300 3468.140 ;
        RECT 2919.700 3465.140 2952.600 3468.140 ;
        RECT -28.380 3465.130 -25.380 3465.140 ;
        RECT 2945.000 3465.130 2948.000 3465.140 ;
        RECT -28.380 3288.140 -25.380 3288.150 ;
        RECT 2945.000 3288.140 2948.000 3288.150 ;
        RECT -32.980 3285.140 0.300 3288.140 ;
        RECT 2919.700 3285.140 2952.600 3288.140 ;
        RECT -28.380 3285.130 -25.380 3285.140 ;
        RECT 2945.000 3285.130 2948.000 3285.140 ;
        RECT -28.380 3108.140 -25.380 3108.150 ;
        RECT 2945.000 3108.140 2948.000 3108.150 ;
        RECT -32.980 3105.140 0.300 3108.140 ;
        RECT 2919.700 3105.140 2952.600 3108.140 ;
        RECT -28.380 3105.130 -25.380 3105.140 ;
        RECT 2945.000 3105.130 2948.000 3105.140 ;
        RECT -28.380 2928.140 -25.380 2928.150 ;
        RECT 2945.000 2928.140 2948.000 2928.150 ;
        RECT -32.980 2925.140 0.300 2928.140 ;
        RECT 2919.700 2925.140 2952.600 2928.140 ;
        RECT -28.380 2925.130 -25.380 2925.140 ;
        RECT 2945.000 2925.130 2948.000 2925.140 ;
        RECT -28.380 2748.140 -25.380 2748.150 ;
        RECT 2945.000 2748.140 2948.000 2748.150 ;
        RECT -32.980 2745.140 0.300 2748.140 ;
        RECT 2919.700 2745.140 2952.600 2748.140 ;
        RECT -28.380 2745.130 -25.380 2745.140 ;
        RECT 2945.000 2745.130 2948.000 2745.140 ;
        RECT -28.380 2568.140 -25.380 2568.150 ;
        RECT 2945.000 2568.140 2948.000 2568.150 ;
        RECT -32.980 2565.140 0.300 2568.140 ;
        RECT 2919.700 2565.140 2952.600 2568.140 ;
        RECT -28.380 2565.130 -25.380 2565.140 ;
        RECT 2945.000 2565.130 2948.000 2565.140 ;
        RECT -28.380 2388.140 -25.380 2388.150 ;
        RECT 2945.000 2388.140 2948.000 2388.150 ;
        RECT -32.980 2385.140 0.300 2388.140 ;
        RECT 2919.700 2385.140 2952.600 2388.140 ;
        RECT -28.380 2385.130 -25.380 2385.140 ;
        RECT 2945.000 2385.130 2948.000 2385.140 ;
        RECT -28.380 2208.140 -25.380 2208.150 ;
        RECT 2945.000 2208.140 2948.000 2208.150 ;
        RECT -32.980 2205.140 0.300 2208.140 ;
        RECT 2919.700 2205.140 2952.600 2208.140 ;
        RECT -28.380 2205.130 -25.380 2205.140 ;
        RECT 2945.000 2205.130 2948.000 2205.140 ;
        RECT -28.380 2028.140 -25.380 2028.150 ;
        RECT 2945.000 2028.140 2948.000 2028.150 ;
        RECT -32.980 2025.140 0.300 2028.140 ;
        RECT 2919.700 2025.140 2952.600 2028.140 ;
        RECT -28.380 2025.130 -25.380 2025.140 ;
        RECT 2945.000 2025.130 2948.000 2025.140 ;
        RECT -28.380 1848.140 -25.380 1848.150 ;
        RECT 2945.000 1848.140 2948.000 1848.150 ;
        RECT -32.980 1845.140 0.300 1848.140 ;
        RECT 2919.700 1845.140 2952.600 1848.140 ;
        RECT -28.380 1845.130 -25.380 1845.140 ;
        RECT 2945.000 1845.130 2948.000 1845.140 ;
        RECT -28.380 1668.140 -25.380 1668.150 ;
        RECT 2945.000 1668.140 2948.000 1668.150 ;
        RECT -32.980 1665.140 0.300 1668.140 ;
        RECT 2919.700 1665.140 2952.600 1668.140 ;
        RECT -28.380 1665.130 -25.380 1665.140 ;
        RECT 2945.000 1665.130 2948.000 1665.140 ;
        RECT -28.380 1488.140 -25.380 1488.150 ;
        RECT 2945.000 1488.140 2948.000 1488.150 ;
        RECT -32.980 1485.140 0.300 1488.140 ;
        RECT 2919.700 1485.140 2952.600 1488.140 ;
        RECT -28.380 1485.130 -25.380 1485.140 ;
        RECT 2945.000 1485.130 2948.000 1485.140 ;
        RECT -28.380 1308.140 -25.380 1308.150 ;
        RECT 2945.000 1308.140 2948.000 1308.150 ;
        RECT -32.980 1305.140 0.300 1308.140 ;
        RECT 2919.700 1305.140 2952.600 1308.140 ;
        RECT -28.380 1305.130 -25.380 1305.140 ;
        RECT 2945.000 1305.130 2948.000 1305.140 ;
        RECT -28.380 1128.140 -25.380 1128.150 ;
        RECT 2945.000 1128.140 2948.000 1128.150 ;
        RECT -32.980 1125.140 0.300 1128.140 ;
        RECT 2919.700 1125.140 2952.600 1128.140 ;
        RECT -28.380 1125.130 -25.380 1125.140 ;
        RECT 2945.000 1125.130 2948.000 1125.140 ;
        RECT -28.380 948.140 -25.380 948.150 ;
        RECT 2945.000 948.140 2948.000 948.150 ;
        RECT -32.980 945.140 0.300 948.140 ;
        RECT 2919.700 945.140 2952.600 948.140 ;
        RECT -28.380 945.130 -25.380 945.140 ;
        RECT 2945.000 945.130 2948.000 945.140 ;
        RECT -28.380 768.140 -25.380 768.150 ;
        RECT 2945.000 768.140 2948.000 768.150 ;
        RECT -32.980 765.140 0.300 768.140 ;
        RECT 2919.700 765.140 2952.600 768.140 ;
        RECT -28.380 765.130 -25.380 765.140 ;
        RECT 2945.000 765.130 2948.000 765.140 ;
        RECT -28.380 588.140 -25.380 588.150 ;
        RECT 2945.000 588.140 2948.000 588.150 ;
        RECT -32.980 585.140 0.300 588.140 ;
        RECT 2919.700 585.140 2952.600 588.140 ;
        RECT -28.380 585.130 -25.380 585.140 ;
        RECT 2945.000 585.130 2948.000 585.140 ;
        RECT -28.380 408.140 -25.380 408.150 ;
        RECT 2945.000 408.140 2948.000 408.150 ;
        RECT -32.980 405.140 0.300 408.140 ;
        RECT 2919.700 405.140 2952.600 408.140 ;
        RECT -28.380 405.130 -25.380 405.140 ;
        RECT 2945.000 405.130 2948.000 405.140 ;
        RECT -28.380 228.140 -25.380 228.150 ;
        RECT 2945.000 228.140 2948.000 228.150 ;
        RECT -32.980 225.140 0.300 228.140 ;
        RECT 2919.700 225.140 2952.600 228.140 ;
        RECT -28.380 225.130 -25.380 225.140 ;
        RECT 2945.000 225.130 2948.000 225.140 ;
        RECT -28.380 48.140 -25.380 48.150 ;
        RECT 2945.000 48.140 2948.000 48.150 ;
        RECT -32.980 45.140 0.300 48.140 ;
        RECT 2919.700 45.140 2952.600 48.140 ;
        RECT -28.380 45.130 -25.380 45.140 ;
        RECT 2945.000 45.130 2948.000 45.140 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 3519.700 133.020 3547.300 ;
        RECT 310.020 3519.700 313.020 3547.300 ;
        RECT 490.020 3519.700 493.020 3547.300 ;
        RECT 670.020 3519.700 673.020 3547.300 ;
        RECT 850.020 3519.700 853.020 3547.300 ;
        RECT 1030.020 3519.700 1033.020 3547.300 ;
        RECT 1210.020 3519.700 1213.020 3547.300 ;
        RECT 1390.020 3519.700 1393.020 3547.300 ;
        RECT 1570.020 3519.700 1573.020 3547.300 ;
        RECT 1750.020 3519.700 1753.020 3547.300 ;
        RECT 1930.020 3519.700 1933.020 3547.300 ;
        RECT 2110.020 3519.700 2113.020 3547.300 ;
        RECT 2290.020 3519.700 2293.020 3547.300 ;
        RECT 2470.020 3519.700 2473.020 3547.300 ;
        RECT 2650.020 3519.700 2653.020 3547.300 ;
        RECT 2830.020 3519.700 2833.020 3547.300 ;
        RECT 130.020 -27.620 133.020 0.300 ;
        RECT 310.020 -27.620 313.020 0.300 ;
        RECT 490.020 -27.620 493.020 0.300 ;
        RECT 670.020 -27.620 673.020 0.300 ;
        RECT 850.020 -27.620 853.020 0.300 ;
        RECT 1030.020 -27.620 1033.020 0.300 ;
        RECT 1210.020 -27.620 1213.020 0.300 ;
        RECT 1390.020 -27.620 1393.020 0.300 ;
        RECT 1570.020 -27.620 1573.020 0.300 ;
        RECT 1750.020 -27.620 1753.020 0.300 ;
        RECT 1930.020 -27.620 1933.020 0.300 ;
        RECT 2110.020 -27.620 2113.020 0.300 ;
        RECT 2290.020 -27.620 2293.020 0.300 ;
        RECT 2470.020 -27.620 2473.020 0.300 ;
        RECT 2650.020 -27.620 2653.020 0.300 ;
        RECT 2830.020 -27.620 2833.020 0.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT -32.070 3376.850 -30.890 3378.030 ;
        RECT -32.070 3375.250 -30.890 3376.430 ;
        RECT -32.070 3196.850 -30.890 3198.030 ;
        RECT -32.070 3195.250 -30.890 3196.430 ;
        RECT -32.070 3016.850 -30.890 3018.030 ;
        RECT -32.070 3015.250 -30.890 3016.430 ;
        RECT -32.070 2836.850 -30.890 2838.030 ;
        RECT -32.070 2835.250 -30.890 2836.430 ;
        RECT -32.070 2656.850 -30.890 2658.030 ;
        RECT -32.070 2655.250 -30.890 2656.430 ;
        RECT -32.070 2476.850 -30.890 2478.030 ;
        RECT -32.070 2475.250 -30.890 2476.430 ;
        RECT -32.070 2296.850 -30.890 2298.030 ;
        RECT -32.070 2295.250 -30.890 2296.430 ;
        RECT -32.070 2116.850 -30.890 2118.030 ;
        RECT -32.070 2115.250 -30.890 2116.430 ;
        RECT -32.070 1936.850 -30.890 1938.030 ;
        RECT -32.070 1935.250 -30.890 1936.430 ;
        RECT -32.070 1756.850 -30.890 1758.030 ;
        RECT -32.070 1755.250 -30.890 1756.430 ;
        RECT -32.070 1576.850 -30.890 1578.030 ;
        RECT -32.070 1575.250 -30.890 1576.430 ;
        RECT -32.070 1396.850 -30.890 1398.030 ;
        RECT -32.070 1395.250 -30.890 1396.430 ;
        RECT -32.070 1216.850 -30.890 1218.030 ;
        RECT -32.070 1215.250 -30.890 1216.430 ;
        RECT -32.070 1036.850 -30.890 1038.030 ;
        RECT -32.070 1035.250 -30.890 1036.430 ;
        RECT -32.070 856.850 -30.890 858.030 ;
        RECT -32.070 855.250 -30.890 856.430 ;
        RECT -32.070 676.850 -30.890 678.030 ;
        RECT -32.070 675.250 -30.890 676.430 ;
        RECT -32.070 496.850 -30.890 498.030 ;
        RECT -32.070 495.250 -30.890 496.430 ;
        RECT -32.070 316.850 -30.890 318.030 ;
        RECT -32.070 315.250 -30.890 316.430 ;
        RECT -32.070 136.850 -30.890 138.030 ;
        RECT -32.070 135.250 -30.890 136.430 ;
        RECT 2950.510 3376.850 2951.690 3378.030 ;
        RECT 2950.510 3375.250 2951.690 3376.430 ;
        RECT 2950.510 3196.850 2951.690 3198.030 ;
        RECT 2950.510 3195.250 2951.690 3196.430 ;
        RECT 2950.510 3016.850 2951.690 3018.030 ;
        RECT 2950.510 3015.250 2951.690 3016.430 ;
        RECT 2950.510 2836.850 2951.690 2838.030 ;
        RECT 2950.510 2835.250 2951.690 2836.430 ;
        RECT 2950.510 2656.850 2951.690 2658.030 ;
        RECT 2950.510 2655.250 2951.690 2656.430 ;
        RECT 2950.510 2476.850 2951.690 2478.030 ;
        RECT 2950.510 2475.250 2951.690 2476.430 ;
        RECT 2950.510 2296.850 2951.690 2298.030 ;
        RECT 2950.510 2295.250 2951.690 2296.430 ;
        RECT 2950.510 2116.850 2951.690 2118.030 ;
        RECT 2950.510 2115.250 2951.690 2116.430 ;
        RECT 2950.510 1936.850 2951.690 1938.030 ;
        RECT 2950.510 1935.250 2951.690 1936.430 ;
        RECT 2950.510 1756.850 2951.690 1758.030 ;
        RECT 2950.510 1755.250 2951.690 1756.430 ;
        RECT 2950.510 1576.850 2951.690 1578.030 ;
        RECT 2950.510 1575.250 2951.690 1576.430 ;
        RECT 2950.510 1396.850 2951.690 1398.030 ;
        RECT 2950.510 1395.250 2951.690 1396.430 ;
        RECT 2950.510 1216.850 2951.690 1218.030 ;
        RECT 2950.510 1215.250 2951.690 1216.430 ;
        RECT 2950.510 1036.850 2951.690 1038.030 ;
        RECT 2950.510 1035.250 2951.690 1036.430 ;
        RECT 2950.510 856.850 2951.690 858.030 ;
        RECT 2950.510 855.250 2951.690 856.430 ;
        RECT 2950.510 676.850 2951.690 678.030 ;
        RECT 2950.510 675.250 2951.690 676.430 ;
        RECT 2950.510 496.850 2951.690 498.030 ;
        RECT 2950.510 495.250 2951.690 496.430 ;
        RECT 2950.510 316.850 2951.690 318.030 ;
        RECT 2950.510 315.250 2951.690 316.430 ;
        RECT 2950.510 136.850 2951.690 138.030 ;
        RECT 2950.510 135.250 2951.690 136.430 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.140 -29.980 3378.150 ;
        RECT 2949.600 3378.140 2952.600 3378.150 ;
        RECT -32.980 3375.140 0.300 3378.140 ;
        RECT 2919.700 3375.140 2952.600 3378.140 ;
        RECT -32.980 3375.130 -29.980 3375.140 ;
        RECT 2949.600 3375.130 2952.600 3375.140 ;
        RECT -32.980 3198.140 -29.980 3198.150 ;
        RECT 2949.600 3198.140 2952.600 3198.150 ;
        RECT -32.980 3195.140 0.300 3198.140 ;
        RECT 2919.700 3195.140 2952.600 3198.140 ;
        RECT -32.980 3195.130 -29.980 3195.140 ;
        RECT 2949.600 3195.130 2952.600 3195.140 ;
        RECT -32.980 3018.140 -29.980 3018.150 ;
        RECT 2949.600 3018.140 2952.600 3018.150 ;
        RECT -32.980 3015.140 0.300 3018.140 ;
        RECT 2919.700 3015.140 2952.600 3018.140 ;
        RECT -32.980 3015.130 -29.980 3015.140 ;
        RECT 2949.600 3015.130 2952.600 3015.140 ;
        RECT -32.980 2838.140 -29.980 2838.150 ;
        RECT 2949.600 2838.140 2952.600 2838.150 ;
        RECT -32.980 2835.140 0.300 2838.140 ;
        RECT 2919.700 2835.140 2952.600 2838.140 ;
        RECT -32.980 2835.130 -29.980 2835.140 ;
        RECT 2949.600 2835.130 2952.600 2835.140 ;
        RECT -32.980 2658.140 -29.980 2658.150 ;
        RECT 2949.600 2658.140 2952.600 2658.150 ;
        RECT -32.980 2655.140 0.300 2658.140 ;
        RECT 2919.700 2655.140 2952.600 2658.140 ;
        RECT -32.980 2655.130 -29.980 2655.140 ;
        RECT 2949.600 2655.130 2952.600 2655.140 ;
        RECT -32.980 2478.140 -29.980 2478.150 ;
        RECT 2949.600 2478.140 2952.600 2478.150 ;
        RECT -32.980 2475.140 0.300 2478.140 ;
        RECT 2919.700 2475.140 2952.600 2478.140 ;
        RECT -32.980 2475.130 -29.980 2475.140 ;
        RECT 2949.600 2475.130 2952.600 2475.140 ;
        RECT -32.980 2298.140 -29.980 2298.150 ;
        RECT 2949.600 2298.140 2952.600 2298.150 ;
        RECT -32.980 2295.140 0.300 2298.140 ;
        RECT 2919.700 2295.140 2952.600 2298.140 ;
        RECT -32.980 2295.130 -29.980 2295.140 ;
        RECT 2949.600 2295.130 2952.600 2295.140 ;
        RECT -32.980 2118.140 -29.980 2118.150 ;
        RECT 2949.600 2118.140 2952.600 2118.150 ;
        RECT -32.980 2115.140 0.300 2118.140 ;
        RECT 2919.700 2115.140 2952.600 2118.140 ;
        RECT -32.980 2115.130 -29.980 2115.140 ;
        RECT 2949.600 2115.130 2952.600 2115.140 ;
        RECT -32.980 1938.140 -29.980 1938.150 ;
        RECT 2949.600 1938.140 2952.600 1938.150 ;
        RECT -32.980 1935.140 0.300 1938.140 ;
        RECT 2919.700 1935.140 2952.600 1938.140 ;
        RECT -32.980 1935.130 -29.980 1935.140 ;
        RECT 2949.600 1935.130 2952.600 1935.140 ;
        RECT -32.980 1758.140 -29.980 1758.150 ;
        RECT 2949.600 1758.140 2952.600 1758.150 ;
        RECT -32.980 1755.140 0.300 1758.140 ;
        RECT 2919.700 1755.140 2952.600 1758.140 ;
        RECT -32.980 1755.130 -29.980 1755.140 ;
        RECT 2949.600 1755.130 2952.600 1755.140 ;
        RECT -32.980 1578.140 -29.980 1578.150 ;
        RECT 2949.600 1578.140 2952.600 1578.150 ;
        RECT -32.980 1575.140 0.300 1578.140 ;
        RECT 2919.700 1575.140 2952.600 1578.140 ;
        RECT -32.980 1575.130 -29.980 1575.140 ;
        RECT 2949.600 1575.130 2952.600 1575.140 ;
        RECT -32.980 1398.140 -29.980 1398.150 ;
        RECT 2949.600 1398.140 2952.600 1398.150 ;
        RECT -32.980 1395.140 0.300 1398.140 ;
        RECT 2919.700 1395.140 2952.600 1398.140 ;
        RECT -32.980 1395.130 -29.980 1395.140 ;
        RECT 2949.600 1395.130 2952.600 1395.140 ;
        RECT -32.980 1218.140 -29.980 1218.150 ;
        RECT 2949.600 1218.140 2952.600 1218.150 ;
        RECT -32.980 1215.140 0.300 1218.140 ;
        RECT 2919.700 1215.140 2952.600 1218.140 ;
        RECT -32.980 1215.130 -29.980 1215.140 ;
        RECT 2949.600 1215.130 2952.600 1215.140 ;
        RECT -32.980 1038.140 -29.980 1038.150 ;
        RECT 2949.600 1038.140 2952.600 1038.150 ;
        RECT -32.980 1035.140 0.300 1038.140 ;
        RECT 2919.700 1035.140 2952.600 1038.140 ;
        RECT -32.980 1035.130 -29.980 1035.140 ;
        RECT 2949.600 1035.130 2952.600 1035.140 ;
        RECT -32.980 858.140 -29.980 858.150 ;
        RECT 2949.600 858.140 2952.600 858.150 ;
        RECT -32.980 855.140 0.300 858.140 ;
        RECT 2919.700 855.140 2952.600 858.140 ;
        RECT -32.980 855.130 -29.980 855.140 ;
        RECT 2949.600 855.130 2952.600 855.140 ;
        RECT -32.980 678.140 -29.980 678.150 ;
        RECT 2949.600 678.140 2952.600 678.150 ;
        RECT -32.980 675.140 0.300 678.140 ;
        RECT 2919.700 675.140 2952.600 678.140 ;
        RECT -32.980 675.130 -29.980 675.140 ;
        RECT 2949.600 675.130 2952.600 675.140 ;
        RECT -32.980 498.140 -29.980 498.150 ;
        RECT 2949.600 498.140 2952.600 498.150 ;
        RECT -32.980 495.140 0.300 498.140 ;
        RECT 2919.700 495.140 2952.600 498.140 ;
        RECT -32.980 495.130 -29.980 495.140 ;
        RECT 2949.600 495.130 2952.600 495.140 ;
        RECT -32.980 318.140 -29.980 318.150 ;
        RECT 2949.600 318.140 2952.600 318.150 ;
        RECT -32.980 315.140 0.300 318.140 ;
        RECT 2919.700 315.140 2952.600 318.140 ;
        RECT -32.980 315.130 -29.980 315.140 ;
        RECT 2949.600 315.130 2952.600 315.140 ;
        RECT -32.980 138.140 -29.980 138.150 ;
        RECT 2949.600 138.140 2952.600 138.150 ;
        RECT -32.980 135.140 0.300 138.140 ;
        RECT 2919.700 135.140 2952.600 138.140 ;
        RECT -32.980 135.130 -29.980 135.140 ;
        RECT 2949.600 135.130 2952.600 135.140 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 3519.700 61.020 3556.500 ;
        RECT 238.020 3519.700 241.020 3556.500 ;
        RECT 418.020 3519.700 421.020 3556.500 ;
        RECT 598.020 3519.700 601.020 3556.500 ;
        RECT 778.020 3519.700 781.020 3556.500 ;
        RECT 958.020 3519.700 961.020 3556.500 ;
        RECT 1138.020 3519.700 1141.020 3556.500 ;
        RECT 1318.020 3519.700 1321.020 3556.500 ;
        RECT 1498.020 3519.700 1501.020 3556.500 ;
        RECT 1678.020 3519.700 1681.020 3556.500 ;
        RECT 1858.020 3519.700 1861.020 3556.500 ;
        RECT 2038.020 3519.700 2041.020 3556.500 ;
        RECT 2218.020 3519.700 2221.020 3556.500 ;
        RECT 2398.020 3519.700 2401.020 3556.500 ;
        RECT 2578.020 3519.700 2581.020 3556.500 ;
        RECT 2758.020 3519.700 2761.020 3556.500 ;
        RECT 58.020 -36.820 61.020 0.300 ;
        RECT 238.020 -36.820 241.020 0.300 ;
        RECT 418.020 -36.820 421.020 0.300 ;
        RECT 598.020 -36.820 601.020 0.300 ;
        RECT 778.020 -36.820 781.020 0.300 ;
        RECT 958.020 -36.820 961.020 0.300 ;
        RECT 1138.020 -36.820 1141.020 0.300 ;
        RECT 1318.020 -36.820 1321.020 0.300 ;
        RECT 1498.020 -36.820 1501.020 0.300 ;
        RECT 1678.020 -36.820 1681.020 0.300 ;
        RECT 1858.020 -36.820 1861.020 0.300 ;
        RECT 2038.020 -36.820 2041.020 0.300 ;
        RECT 2218.020 -36.820 2221.020 0.300 ;
        RECT 2398.020 -36.820 2401.020 0.300 ;
        RECT 2578.020 -36.820 2581.020 0.300 ;
        RECT 2758.020 -36.820 2761.020 0.300 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT -36.670 3484.850 -35.490 3486.030 ;
        RECT -36.670 3483.250 -35.490 3484.430 ;
        RECT -36.670 3304.850 -35.490 3306.030 ;
        RECT -36.670 3303.250 -35.490 3304.430 ;
        RECT -36.670 3124.850 -35.490 3126.030 ;
        RECT -36.670 3123.250 -35.490 3124.430 ;
        RECT -36.670 2944.850 -35.490 2946.030 ;
        RECT -36.670 2943.250 -35.490 2944.430 ;
        RECT -36.670 2764.850 -35.490 2766.030 ;
        RECT -36.670 2763.250 -35.490 2764.430 ;
        RECT -36.670 2584.850 -35.490 2586.030 ;
        RECT -36.670 2583.250 -35.490 2584.430 ;
        RECT -36.670 2404.850 -35.490 2406.030 ;
        RECT -36.670 2403.250 -35.490 2404.430 ;
        RECT -36.670 2224.850 -35.490 2226.030 ;
        RECT -36.670 2223.250 -35.490 2224.430 ;
        RECT -36.670 2044.850 -35.490 2046.030 ;
        RECT -36.670 2043.250 -35.490 2044.430 ;
        RECT -36.670 1864.850 -35.490 1866.030 ;
        RECT -36.670 1863.250 -35.490 1864.430 ;
        RECT -36.670 1684.850 -35.490 1686.030 ;
        RECT -36.670 1683.250 -35.490 1684.430 ;
        RECT -36.670 1504.850 -35.490 1506.030 ;
        RECT -36.670 1503.250 -35.490 1504.430 ;
        RECT -36.670 1324.850 -35.490 1326.030 ;
        RECT -36.670 1323.250 -35.490 1324.430 ;
        RECT -36.670 1144.850 -35.490 1146.030 ;
        RECT -36.670 1143.250 -35.490 1144.430 ;
        RECT -36.670 964.850 -35.490 966.030 ;
        RECT -36.670 963.250 -35.490 964.430 ;
        RECT -36.670 784.850 -35.490 786.030 ;
        RECT -36.670 783.250 -35.490 784.430 ;
        RECT -36.670 604.850 -35.490 606.030 ;
        RECT -36.670 603.250 -35.490 604.430 ;
        RECT -36.670 424.850 -35.490 426.030 ;
        RECT -36.670 423.250 -35.490 424.430 ;
        RECT -36.670 244.850 -35.490 246.030 ;
        RECT -36.670 243.250 -35.490 244.430 ;
        RECT -36.670 64.850 -35.490 66.030 ;
        RECT -36.670 63.250 -35.490 64.430 ;
        RECT 2955.110 3484.850 2956.290 3486.030 ;
        RECT 2955.110 3483.250 2956.290 3484.430 ;
        RECT 2955.110 3304.850 2956.290 3306.030 ;
        RECT 2955.110 3303.250 2956.290 3304.430 ;
        RECT 2955.110 3124.850 2956.290 3126.030 ;
        RECT 2955.110 3123.250 2956.290 3124.430 ;
        RECT 2955.110 2944.850 2956.290 2946.030 ;
        RECT 2955.110 2943.250 2956.290 2944.430 ;
        RECT 2955.110 2764.850 2956.290 2766.030 ;
        RECT 2955.110 2763.250 2956.290 2764.430 ;
        RECT 2955.110 2584.850 2956.290 2586.030 ;
        RECT 2955.110 2583.250 2956.290 2584.430 ;
        RECT 2955.110 2404.850 2956.290 2406.030 ;
        RECT 2955.110 2403.250 2956.290 2404.430 ;
        RECT 2955.110 2224.850 2956.290 2226.030 ;
        RECT 2955.110 2223.250 2956.290 2224.430 ;
        RECT 2955.110 2044.850 2956.290 2046.030 ;
        RECT 2955.110 2043.250 2956.290 2044.430 ;
        RECT 2955.110 1864.850 2956.290 1866.030 ;
        RECT 2955.110 1863.250 2956.290 1864.430 ;
        RECT 2955.110 1684.850 2956.290 1686.030 ;
        RECT 2955.110 1683.250 2956.290 1684.430 ;
        RECT 2955.110 1504.850 2956.290 1506.030 ;
        RECT 2955.110 1503.250 2956.290 1504.430 ;
        RECT 2955.110 1324.850 2956.290 1326.030 ;
        RECT 2955.110 1323.250 2956.290 1324.430 ;
        RECT 2955.110 1144.850 2956.290 1146.030 ;
        RECT 2955.110 1143.250 2956.290 1144.430 ;
        RECT 2955.110 964.850 2956.290 966.030 ;
        RECT 2955.110 963.250 2956.290 964.430 ;
        RECT 2955.110 784.850 2956.290 786.030 ;
        RECT 2955.110 783.250 2956.290 784.430 ;
        RECT 2955.110 604.850 2956.290 606.030 ;
        RECT 2955.110 603.250 2956.290 604.430 ;
        RECT 2955.110 424.850 2956.290 426.030 ;
        RECT 2955.110 423.250 2956.290 424.430 ;
        RECT 2955.110 244.850 2956.290 246.030 ;
        RECT 2955.110 243.250 2956.290 244.430 ;
        RECT 2955.110 64.850 2956.290 66.030 ;
        RECT 2955.110 63.250 2956.290 64.430 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.140 -34.580 3486.150 ;
        RECT 2954.200 3486.140 2957.200 3486.150 ;
        RECT -42.180 3483.140 0.300 3486.140 ;
        RECT 2919.700 3483.140 2961.800 3486.140 ;
        RECT -37.580 3483.130 -34.580 3483.140 ;
        RECT 2954.200 3483.130 2957.200 3483.140 ;
        RECT -37.580 3306.140 -34.580 3306.150 ;
        RECT 2954.200 3306.140 2957.200 3306.150 ;
        RECT -42.180 3303.140 0.300 3306.140 ;
        RECT 2919.700 3303.140 2961.800 3306.140 ;
        RECT -37.580 3303.130 -34.580 3303.140 ;
        RECT 2954.200 3303.130 2957.200 3303.140 ;
        RECT -37.580 3126.140 -34.580 3126.150 ;
        RECT 2954.200 3126.140 2957.200 3126.150 ;
        RECT -42.180 3123.140 0.300 3126.140 ;
        RECT 2919.700 3123.140 2961.800 3126.140 ;
        RECT -37.580 3123.130 -34.580 3123.140 ;
        RECT 2954.200 3123.130 2957.200 3123.140 ;
        RECT -37.580 2946.140 -34.580 2946.150 ;
        RECT 2954.200 2946.140 2957.200 2946.150 ;
        RECT -42.180 2943.140 0.300 2946.140 ;
        RECT 2919.700 2943.140 2961.800 2946.140 ;
        RECT -37.580 2943.130 -34.580 2943.140 ;
        RECT 2954.200 2943.130 2957.200 2943.140 ;
        RECT -37.580 2766.140 -34.580 2766.150 ;
        RECT 2954.200 2766.140 2957.200 2766.150 ;
        RECT -42.180 2763.140 0.300 2766.140 ;
        RECT 2919.700 2763.140 2961.800 2766.140 ;
        RECT -37.580 2763.130 -34.580 2763.140 ;
        RECT 2954.200 2763.130 2957.200 2763.140 ;
        RECT -37.580 2586.140 -34.580 2586.150 ;
        RECT 2954.200 2586.140 2957.200 2586.150 ;
        RECT -42.180 2583.140 0.300 2586.140 ;
        RECT 2919.700 2583.140 2961.800 2586.140 ;
        RECT -37.580 2583.130 -34.580 2583.140 ;
        RECT 2954.200 2583.130 2957.200 2583.140 ;
        RECT -37.580 2406.140 -34.580 2406.150 ;
        RECT 2954.200 2406.140 2957.200 2406.150 ;
        RECT -42.180 2403.140 0.300 2406.140 ;
        RECT 2919.700 2403.140 2961.800 2406.140 ;
        RECT -37.580 2403.130 -34.580 2403.140 ;
        RECT 2954.200 2403.130 2957.200 2403.140 ;
        RECT -37.580 2226.140 -34.580 2226.150 ;
        RECT 2954.200 2226.140 2957.200 2226.150 ;
        RECT -42.180 2223.140 0.300 2226.140 ;
        RECT 2919.700 2223.140 2961.800 2226.140 ;
        RECT -37.580 2223.130 -34.580 2223.140 ;
        RECT 2954.200 2223.130 2957.200 2223.140 ;
        RECT -37.580 2046.140 -34.580 2046.150 ;
        RECT 2954.200 2046.140 2957.200 2046.150 ;
        RECT -42.180 2043.140 0.300 2046.140 ;
        RECT 2919.700 2043.140 2961.800 2046.140 ;
        RECT -37.580 2043.130 -34.580 2043.140 ;
        RECT 2954.200 2043.130 2957.200 2043.140 ;
        RECT -37.580 1866.140 -34.580 1866.150 ;
        RECT 2954.200 1866.140 2957.200 1866.150 ;
        RECT -42.180 1863.140 0.300 1866.140 ;
        RECT 2919.700 1863.140 2961.800 1866.140 ;
        RECT -37.580 1863.130 -34.580 1863.140 ;
        RECT 2954.200 1863.130 2957.200 1863.140 ;
        RECT -37.580 1686.140 -34.580 1686.150 ;
        RECT 2954.200 1686.140 2957.200 1686.150 ;
        RECT -42.180 1683.140 0.300 1686.140 ;
        RECT 2919.700 1683.140 2961.800 1686.140 ;
        RECT -37.580 1683.130 -34.580 1683.140 ;
        RECT 2954.200 1683.130 2957.200 1683.140 ;
        RECT -37.580 1506.140 -34.580 1506.150 ;
        RECT 2954.200 1506.140 2957.200 1506.150 ;
        RECT -42.180 1503.140 0.300 1506.140 ;
        RECT 2919.700 1503.140 2961.800 1506.140 ;
        RECT -37.580 1503.130 -34.580 1503.140 ;
        RECT 2954.200 1503.130 2957.200 1503.140 ;
        RECT -37.580 1326.140 -34.580 1326.150 ;
        RECT 2954.200 1326.140 2957.200 1326.150 ;
        RECT -42.180 1323.140 0.300 1326.140 ;
        RECT 2919.700 1323.140 2961.800 1326.140 ;
        RECT -37.580 1323.130 -34.580 1323.140 ;
        RECT 2954.200 1323.130 2957.200 1323.140 ;
        RECT -37.580 1146.140 -34.580 1146.150 ;
        RECT 2954.200 1146.140 2957.200 1146.150 ;
        RECT -42.180 1143.140 0.300 1146.140 ;
        RECT 2919.700 1143.140 2961.800 1146.140 ;
        RECT -37.580 1143.130 -34.580 1143.140 ;
        RECT 2954.200 1143.130 2957.200 1143.140 ;
        RECT -37.580 966.140 -34.580 966.150 ;
        RECT 2954.200 966.140 2957.200 966.150 ;
        RECT -42.180 963.140 0.300 966.140 ;
        RECT 2919.700 963.140 2961.800 966.140 ;
        RECT -37.580 963.130 -34.580 963.140 ;
        RECT 2954.200 963.130 2957.200 963.140 ;
        RECT -37.580 786.140 -34.580 786.150 ;
        RECT 2954.200 786.140 2957.200 786.150 ;
        RECT -42.180 783.140 0.300 786.140 ;
        RECT 2919.700 783.140 2961.800 786.140 ;
        RECT -37.580 783.130 -34.580 783.140 ;
        RECT 2954.200 783.130 2957.200 783.140 ;
        RECT -37.580 606.140 -34.580 606.150 ;
        RECT 2954.200 606.140 2957.200 606.150 ;
        RECT -42.180 603.140 0.300 606.140 ;
        RECT 2919.700 603.140 2961.800 606.140 ;
        RECT -37.580 603.130 -34.580 603.140 ;
        RECT 2954.200 603.130 2957.200 603.140 ;
        RECT -37.580 426.140 -34.580 426.150 ;
        RECT 2954.200 426.140 2957.200 426.150 ;
        RECT -42.180 423.140 0.300 426.140 ;
        RECT 2919.700 423.140 2961.800 426.140 ;
        RECT -37.580 423.130 -34.580 423.140 ;
        RECT 2954.200 423.130 2957.200 423.140 ;
        RECT -37.580 246.140 -34.580 246.150 ;
        RECT 2954.200 246.140 2957.200 246.150 ;
        RECT -42.180 243.140 0.300 246.140 ;
        RECT 2919.700 243.140 2961.800 246.140 ;
        RECT -37.580 243.130 -34.580 243.140 ;
        RECT 2954.200 243.130 2957.200 243.140 ;
        RECT -37.580 66.140 -34.580 66.150 ;
        RECT 2954.200 66.140 2957.200 66.150 ;
        RECT -42.180 63.140 0.300 66.140 ;
        RECT 2919.700 63.140 2961.800 66.140 ;
        RECT -37.580 63.130 -34.580 63.140 ;
        RECT 2954.200 63.130 2957.200 63.140 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 3519.700 151.020 3556.500 ;
        RECT 328.020 3519.700 331.020 3556.500 ;
        RECT 508.020 3519.700 511.020 3556.500 ;
        RECT 688.020 3519.700 691.020 3556.500 ;
        RECT 868.020 3519.700 871.020 3556.500 ;
        RECT 1048.020 3519.700 1051.020 3556.500 ;
        RECT 1228.020 3519.700 1231.020 3556.500 ;
        RECT 1408.020 3519.700 1411.020 3556.500 ;
        RECT 1588.020 3519.700 1591.020 3556.500 ;
        RECT 1768.020 3519.700 1771.020 3556.500 ;
        RECT 1948.020 3519.700 1951.020 3556.500 ;
        RECT 2128.020 3519.700 2131.020 3556.500 ;
        RECT 2308.020 3519.700 2311.020 3556.500 ;
        RECT 2488.020 3519.700 2491.020 3556.500 ;
        RECT 2668.020 3519.700 2671.020 3556.500 ;
        RECT 2848.020 3519.700 2851.020 3556.500 ;
        RECT 148.020 -36.820 151.020 0.300 ;
        RECT 328.020 -36.820 331.020 0.300 ;
        RECT 508.020 -36.820 511.020 0.300 ;
        RECT 688.020 -36.820 691.020 0.300 ;
        RECT 868.020 -36.820 871.020 0.300 ;
        RECT 1048.020 -36.820 1051.020 0.300 ;
        RECT 1228.020 -36.820 1231.020 0.300 ;
        RECT 1408.020 -36.820 1411.020 0.300 ;
        RECT 1588.020 -36.820 1591.020 0.300 ;
        RECT 1768.020 -36.820 1771.020 0.300 ;
        RECT 1948.020 -36.820 1951.020 0.300 ;
        RECT 2128.020 -36.820 2131.020 0.300 ;
        RECT 2308.020 -36.820 2311.020 0.300 ;
        RECT 2488.020 -36.820 2491.020 0.300 ;
        RECT 2668.020 -36.820 2671.020 0.300 ;
        RECT 2848.020 -36.820 2851.020 0.300 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT -41.270 3394.850 -40.090 3396.030 ;
        RECT -41.270 3393.250 -40.090 3394.430 ;
        RECT -41.270 3214.850 -40.090 3216.030 ;
        RECT -41.270 3213.250 -40.090 3214.430 ;
        RECT -41.270 3034.850 -40.090 3036.030 ;
        RECT -41.270 3033.250 -40.090 3034.430 ;
        RECT -41.270 2854.850 -40.090 2856.030 ;
        RECT -41.270 2853.250 -40.090 2854.430 ;
        RECT -41.270 2674.850 -40.090 2676.030 ;
        RECT -41.270 2673.250 -40.090 2674.430 ;
        RECT -41.270 2494.850 -40.090 2496.030 ;
        RECT -41.270 2493.250 -40.090 2494.430 ;
        RECT -41.270 2314.850 -40.090 2316.030 ;
        RECT -41.270 2313.250 -40.090 2314.430 ;
        RECT -41.270 2134.850 -40.090 2136.030 ;
        RECT -41.270 2133.250 -40.090 2134.430 ;
        RECT -41.270 1954.850 -40.090 1956.030 ;
        RECT -41.270 1953.250 -40.090 1954.430 ;
        RECT -41.270 1774.850 -40.090 1776.030 ;
        RECT -41.270 1773.250 -40.090 1774.430 ;
        RECT -41.270 1594.850 -40.090 1596.030 ;
        RECT -41.270 1593.250 -40.090 1594.430 ;
        RECT -41.270 1414.850 -40.090 1416.030 ;
        RECT -41.270 1413.250 -40.090 1414.430 ;
        RECT -41.270 1234.850 -40.090 1236.030 ;
        RECT -41.270 1233.250 -40.090 1234.430 ;
        RECT -41.270 1054.850 -40.090 1056.030 ;
        RECT -41.270 1053.250 -40.090 1054.430 ;
        RECT -41.270 874.850 -40.090 876.030 ;
        RECT -41.270 873.250 -40.090 874.430 ;
        RECT -41.270 694.850 -40.090 696.030 ;
        RECT -41.270 693.250 -40.090 694.430 ;
        RECT -41.270 514.850 -40.090 516.030 ;
        RECT -41.270 513.250 -40.090 514.430 ;
        RECT -41.270 334.850 -40.090 336.030 ;
        RECT -41.270 333.250 -40.090 334.430 ;
        RECT -41.270 154.850 -40.090 156.030 ;
        RECT -41.270 153.250 -40.090 154.430 ;
        RECT 2959.710 3394.850 2960.890 3396.030 ;
        RECT 2959.710 3393.250 2960.890 3394.430 ;
        RECT 2959.710 3214.850 2960.890 3216.030 ;
        RECT 2959.710 3213.250 2960.890 3214.430 ;
        RECT 2959.710 3034.850 2960.890 3036.030 ;
        RECT 2959.710 3033.250 2960.890 3034.430 ;
        RECT 2959.710 2854.850 2960.890 2856.030 ;
        RECT 2959.710 2853.250 2960.890 2854.430 ;
        RECT 2959.710 2674.850 2960.890 2676.030 ;
        RECT 2959.710 2673.250 2960.890 2674.430 ;
        RECT 2959.710 2494.850 2960.890 2496.030 ;
        RECT 2959.710 2493.250 2960.890 2494.430 ;
        RECT 2959.710 2314.850 2960.890 2316.030 ;
        RECT 2959.710 2313.250 2960.890 2314.430 ;
        RECT 2959.710 2134.850 2960.890 2136.030 ;
        RECT 2959.710 2133.250 2960.890 2134.430 ;
        RECT 2959.710 1954.850 2960.890 1956.030 ;
        RECT 2959.710 1953.250 2960.890 1954.430 ;
        RECT 2959.710 1774.850 2960.890 1776.030 ;
        RECT 2959.710 1773.250 2960.890 1774.430 ;
        RECT 2959.710 1594.850 2960.890 1596.030 ;
        RECT 2959.710 1593.250 2960.890 1594.430 ;
        RECT 2959.710 1414.850 2960.890 1416.030 ;
        RECT 2959.710 1413.250 2960.890 1414.430 ;
        RECT 2959.710 1234.850 2960.890 1236.030 ;
        RECT 2959.710 1233.250 2960.890 1234.430 ;
        RECT 2959.710 1054.850 2960.890 1056.030 ;
        RECT 2959.710 1053.250 2960.890 1054.430 ;
        RECT 2959.710 874.850 2960.890 876.030 ;
        RECT 2959.710 873.250 2960.890 874.430 ;
        RECT 2959.710 694.850 2960.890 696.030 ;
        RECT 2959.710 693.250 2960.890 694.430 ;
        RECT 2959.710 514.850 2960.890 516.030 ;
        RECT 2959.710 513.250 2960.890 514.430 ;
        RECT 2959.710 334.850 2960.890 336.030 ;
        RECT 2959.710 333.250 2960.890 334.430 ;
        RECT 2959.710 154.850 2960.890 156.030 ;
        RECT 2959.710 153.250 2960.890 154.430 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.140 -39.180 3396.150 ;
        RECT 2958.800 3396.140 2961.800 3396.150 ;
        RECT -42.180 3393.140 0.300 3396.140 ;
        RECT 2919.700 3393.140 2961.800 3396.140 ;
        RECT -42.180 3393.130 -39.180 3393.140 ;
        RECT 2958.800 3393.130 2961.800 3393.140 ;
        RECT -42.180 3216.140 -39.180 3216.150 ;
        RECT 2958.800 3216.140 2961.800 3216.150 ;
        RECT -42.180 3213.140 0.300 3216.140 ;
        RECT 2919.700 3213.140 2961.800 3216.140 ;
        RECT -42.180 3213.130 -39.180 3213.140 ;
        RECT 2958.800 3213.130 2961.800 3213.140 ;
        RECT -42.180 3036.140 -39.180 3036.150 ;
        RECT 2958.800 3036.140 2961.800 3036.150 ;
        RECT -42.180 3033.140 0.300 3036.140 ;
        RECT 2919.700 3033.140 2961.800 3036.140 ;
        RECT -42.180 3033.130 -39.180 3033.140 ;
        RECT 2958.800 3033.130 2961.800 3033.140 ;
        RECT -42.180 2856.140 -39.180 2856.150 ;
        RECT 2958.800 2856.140 2961.800 2856.150 ;
        RECT -42.180 2853.140 0.300 2856.140 ;
        RECT 2919.700 2853.140 2961.800 2856.140 ;
        RECT -42.180 2853.130 -39.180 2853.140 ;
        RECT 2958.800 2853.130 2961.800 2853.140 ;
        RECT -42.180 2676.140 -39.180 2676.150 ;
        RECT 2958.800 2676.140 2961.800 2676.150 ;
        RECT -42.180 2673.140 0.300 2676.140 ;
        RECT 2919.700 2673.140 2961.800 2676.140 ;
        RECT -42.180 2673.130 -39.180 2673.140 ;
        RECT 2958.800 2673.130 2961.800 2673.140 ;
        RECT -42.180 2496.140 -39.180 2496.150 ;
        RECT 2958.800 2496.140 2961.800 2496.150 ;
        RECT -42.180 2493.140 0.300 2496.140 ;
        RECT 2919.700 2493.140 2961.800 2496.140 ;
        RECT -42.180 2493.130 -39.180 2493.140 ;
        RECT 2958.800 2493.130 2961.800 2493.140 ;
        RECT -42.180 2316.140 -39.180 2316.150 ;
        RECT 2958.800 2316.140 2961.800 2316.150 ;
        RECT -42.180 2313.140 0.300 2316.140 ;
        RECT 2919.700 2313.140 2961.800 2316.140 ;
        RECT -42.180 2313.130 -39.180 2313.140 ;
        RECT 2958.800 2313.130 2961.800 2313.140 ;
        RECT -42.180 2136.140 -39.180 2136.150 ;
        RECT 2958.800 2136.140 2961.800 2136.150 ;
        RECT -42.180 2133.140 0.300 2136.140 ;
        RECT 2919.700 2133.140 2961.800 2136.140 ;
        RECT -42.180 2133.130 -39.180 2133.140 ;
        RECT 2958.800 2133.130 2961.800 2133.140 ;
        RECT -42.180 1956.140 -39.180 1956.150 ;
        RECT 2958.800 1956.140 2961.800 1956.150 ;
        RECT -42.180 1953.140 0.300 1956.140 ;
        RECT 2919.700 1953.140 2961.800 1956.140 ;
        RECT -42.180 1953.130 -39.180 1953.140 ;
        RECT 2958.800 1953.130 2961.800 1953.140 ;
        RECT -42.180 1776.140 -39.180 1776.150 ;
        RECT 2958.800 1776.140 2961.800 1776.150 ;
        RECT -42.180 1773.140 0.300 1776.140 ;
        RECT 2919.700 1773.140 2961.800 1776.140 ;
        RECT -42.180 1773.130 -39.180 1773.140 ;
        RECT 2958.800 1773.130 2961.800 1773.140 ;
        RECT -42.180 1596.140 -39.180 1596.150 ;
        RECT 2958.800 1596.140 2961.800 1596.150 ;
        RECT -42.180 1593.140 0.300 1596.140 ;
        RECT 2919.700 1593.140 2961.800 1596.140 ;
        RECT -42.180 1593.130 -39.180 1593.140 ;
        RECT 2958.800 1593.130 2961.800 1593.140 ;
        RECT -42.180 1416.140 -39.180 1416.150 ;
        RECT 2958.800 1416.140 2961.800 1416.150 ;
        RECT -42.180 1413.140 0.300 1416.140 ;
        RECT 2919.700 1413.140 2961.800 1416.140 ;
        RECT -42.180 1413.130 -39.180 1413.140 ;
        RECT 2958.800 1413.130 2961.800 1413.140 ;
        RECT -42.180 1236.140 -39.180 1236.150 ;
        RECT 2958.800 1236.140 2961.800 1236.150 ;
        RECT -42.180 1233.140 0.300 1236.140 ;
        RECT 2919.700 1233.140 2961.800 1236.140 ;
        RECT -42.180 1233.130 -39.180 1233.140 ;
        RECT 2958.800 1233.130 2961.800 1233.140 ;
        RECT -42.180 1056.140 -39.180 1056.150 ;
        RECT 2958.800 1056.140 2961.800 1056.150 ;
        RECT -42.180 1053.140 0.300 1056.140 ;
        RECT 2919.700 1053.140 2961.800 1056.140 ;
        RECT -42.180 1053.130 -39.180 1053.140 ;
        RECT 2958.800 1053.130 2961.800 1053.140 ;
        RECT -42.180 876.140 -39.180 876.150 ;
        RECT 2958.800 876.140 2961.800 876.150 ;
        RECT -42.180 873.140 0.300 876.140 ;
        RECT 2919.700 873.140 2961.800 876.140 ;
        RECT -42.180 873.130 -39.180 873.140 ;
        RECT 2958.800 873.130 2961.800 873.140 ;
        RECT -42.180 696.140 -39.180 696.150 ;
        RECT 2958.800 696.140 2961.800 696.150 ;
        RECT -42.180 693.140 0.300 696.140 ;
        RECT 2919.700 693.140 2961.800 696.140 ;
        RECT -42.180 693.130 -39.180 693.140 ;
        RECT 2958.800 693.130 2961.800 693.140 ;
        RECT -42.180 516.140 -39.180 516.150 ;
        RECT 2958.800 516.140 2961.800 516.150 ;
        RECT -42.180 513.140 0.300 516.140 ;
        RECT 2919.700 513.140 2961.800 516.140 ;
        RECT -42.180 513.130 -39.180 513.140 ;
        RECT 2958.800 513.130 2961.800 513.140 ;
        RECT -42.180 336.140 -39.180 336.150 ;
        RECT 2958.800 336.140 2961.800 336.150 ;
        RECT -42.180 333.140 0.300 336.140 ;
        RECT 2919.700 333.140 2961.800 336.140 ;
        RECT -42.180 333.130 -39.180 333.140 ;
        RECT 2958.800 333.130 2961.800 333.140 ;
        RECT -42.180 156.140 -39.180 156.150 ;
        RECT 2958.800 156.140 2961.800 156.150 ;
        RECT -42.180 153.140 0.300 156.140 ;
        RECT 2919.700 153.140 2961.800 156.140 ;
        RECT -42.180 153.130 -39.180 153.140 ;
        RECT 2958.800 153.130 2961.800 153.140 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2914.100 3508.885 ;
      LAYER met1 ;
        RECT 2.830 2.760 2914.100 3509.040 ;
      LAYER met2 ;
        RECT 2.710 0.300 2917.370 3519.700 ;
      LAYER met3 ;
        RECT 0.300 10.715 2919.700 3508.965 ;
      LAYER met4 ;
        RECT 4.020 0.300 2910.090 3519.700 ;
      LAYER met5 ;
        RECT 0.300 9.130 2919.700 3486.140 ;
  END
END user_project_wrapper
END LIBRARY

